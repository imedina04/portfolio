`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mXW6bUl5enO4TRMKolk/ZdGy0k/Wa3ixEOJFdKNe3zr2aDiWN/6uzpH1bLXDjbjJiQ/H/8Zk0tUc
zHB5+a9AOw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YrV3De7K+YpadhprwHFki3u1JYgILJAIDHx8JyzOZ5ZyZe1xsfzrZlhZgo9y1THWLYJVYvRLjLUF
8UECtWGTS9LCbRO6LpIO0zdxMZel9X/wF9NYGduH0LdFZdGHWV20c66Lx1Dmu99WHTe+6bwqgyuK
a5HhHw6Xh2bef5pyVpw=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
r45Vmg2hm2GZWhRHiz3jT8i2aHCx1CpyYm289L9dvMzYfnwa19f39tCi3RwZ1fGScagNb/k8Wvxo
CcTC+NrFMBfIBBz4MvqyZ8IdKL3NAEkUm5koxVgdwyIdDNVYZinySunBz3VWNdsQMi/UdLMIRrky
BoIuydnIik4maDPVlqT4rPCbZpaD1MiTm0V1YtDT89f+NvlGejBWcgOoJ4+oJ927SvJCCSA/2o4L
xIsDpnhNGOzXwq4cNzvcv1Bv6+ImH9ElqfHk5PU843hmKFWaoUJ+XwDBSEllq8FiFhVOdacW+0L3
onLX/ovKi1vmSTrXoYGiH93PU127c8zS/YIuhw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KkNAK9QAtT6wOxT5+WTYnMXJulhUXr5f64M/aLgOG/uGlUv+e6+Tg8Tq3TxUtvqXTbFTAAFbvNwa
A26K0bI4rJ/VHL5cpusuetQlfQQrfNPL+85zGQtFZbIqlPDBG9PvZcgfGkQexKIi1ZIzqEd7J9ae
DjIazpffXnoSf1HprxEPwKGs2CHymtf8zv8RrTiTXwwI1xS1x5MdP927yfx/W3+Dru0teV+3f9vc
iy6q1Bxj6FhygH+4mh2/h7BBuNfeQRQk039twHs/GZ5/MoIqUk/pgsCXLCbq8MF3wtzOteW5DoXr
hpmW54ZRIVFUIUo/Iaf7rXAkjybd2xt1Hbibkg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TEKg+63TKYP3Gmaz+p89Z3UTu5p3NxyuACVHbARoRLL0R77dfUa1QDMfgNuFKg8hIaZLVRsSr/jT
F621qiv1nBzTmeRsKOvSnTksLEnvxgiRZCEOvbU7X/9gCXCZK0B9i4oy4ACYoT6Hq6BvHOL5TI2W
CoFIcCFutl2KPyMXhSace/hSDm4EtiJAQLRpq8XgMGXwRpZ/xdG2Na+BN9vXVHtjY2Vg3npqR5fH
bcNYc0J0HA+9H4BqQ2vphaIfuxV5aMxK5mUwmtLZKYZ5u29ilEBzi/GAN8J59cN3H+8RjJ76r0A3
KhOJ0C+M+z5+Zbw24Vzd/m3p7iiVTp+acnwwxQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XrwB0OVtkmQgH3kKxB3Mo8alTC9ZT2gdavhm/rF7EOnBFqpHvafG2e0WDVO4u/WnticaCcVkYY4B
IlmkwmbTXf2+U151n8NYIhEHoNtbA91rvoWEQ/jPb7rY+1uF9dkLLzaJAr60PuQXXSTBvjnmCV/1
39OIjjSZO6cVv7bDxLA=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AwuPeyMqg/J6Z+iq2u6vpWGK9asqvIBRvw+7fjvyFL64PnhUKzAaSeWYgULuDTuG1QCJwC8+1tM6
vE1UlEAL6iE4hEdSDoDOn6/s2zKYeNu3st3cKLxbB5YZtbXLMTA128F13D5a6y//ApmTjddUjem0
09ihCTQt0jfeDKjmR+m2wMbQrTW/uX4s1hUWCLZ6DIUl6HqUGKJ0Zx/SafYizGEZhm7+AMKrMNLr
ch37HgKjex/XwrEX7qBDlbA5HULUvY1qU7382PUKrvMaRWGodtSD0H+Gtv4pUSI2rlE8IF5i3CiU
H8r7QIWCO1PF40B8fBNDHBgkmitB9zMLWMfWmg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 137008)
`protect data_block
Gtr34gEEe7LAlmRaU77+BpYYw9iOpFAjz2nJzKEnLW+JDq9ObKTbzNKfL4vWz7tR2UzOYXUO1GRn
S/dy0ejutATRGvMaWcSVsB+LdD4oHfa/kkEkk8lg1dfk00clOM2mcPF+Yyyu6g5FgMi0/JN/xxCK
UGU3qhPNv48jZuOee5h2KvT2/NNnOH72Xy9WuAm0IjyU2grLOl60TvKACmYuN3G/IImcVVeibn0l
7Jc88bT6/HY427Roy3U1+qFp/MsDsaw7FAL4QcvEVKtk4IfU7yeyKDOOdrSFWEvM9xLuFJ4eFbTr
Pjyxtq2qtVTQtHPq4v2yJkULntw5UMIB9S8krCshz1cGj7ZW0N2SLDer/s6i091QL8oRPdkvU+4i
UF7on5WKntpn+L5H9nCEs0PyAnhKICb4Chdz7NV1RIHdI/8svIle9z2u+Hqpj0QS8UsetGEAcxh/
Ghg/906pTTlRMsMjedrrXG+tMacD3jd1KE7sLmx5M1DisN6eSgpaQ5+J6ywys9Q6Bz7i+citcxlv
X5F/FR23Bwr5c6fdVf6at1KEc74MPsMbBSbXMBBnJJQZyysPHe4Xu3kkgLgsRT+4FPeLeaX1bmiz
xYme0HxOCi4nVl0iopT9Zlcxh8u2El+lQbmw1uowKPCN8uAVJuWLy/bhLQjq2m8Tu/Bi48yXQz0r
a0nNu/fKp5tggPDs9fqiYLl4Z0i9iy/LMpTjmmkwh8hQ/ah6LJGyKoMFeBbV/G+pcIYlBoDjwSNU
i8iqXuyYrI4k3pqgYksFIvERfkPk8dhCs8a4WbY5k0IaY4odJChsZNaRHgD53bqZoZR/LhZQOQrr
ZDVcMk0rMpG6LwKObG9aMcGIC+i4rPAjNdJiMm0lgG+/hzzXZFHeF0/sS4JXvIr6Hr8AqT+lJkyP
8KxcJ4dapgtzz3uCnloc7fxDA3B8V0SweA/G87sA/TPgOwnjoYHVsySU/rH1GlnwJCoO/5Ve1tzw
fy3JUyc8zudHxTzYG1HZU65gVnDcpdOjOqdSr9WW02f+7qboPGh+FBBOFF+rtG6CaIdj4J3Ejmdo
AVbvymF9dg04fN65OAxz9Qxnhxzap+71/J4vBgntc2lBixu43nUq5vAtEsBTF1jJJAx3zyttW3L0
potsY9IEyZk95vyU6S3YzjAeaPdVvKJftxJnrh1i64yipiHiTBSy0OStdL2gOXxz08jYVUKeAAuV
N1ByhF3M8qgeD7DwPwf2KVv4ieyjbATY6IlAOvykEGLYdkqwzNRCNWCrWILFfEFJ7QNMNREjRBpp
dAqfcBO+bYTbRjr6j+23mMavWugoYFSlLaV1mGOpzSfYIDJvzldn9d+ZzSDA7JQPze1Z3bvYvXl/
CW4gviGJN923sdT60YOkqX1CvcHwM3siYAjWmqijsMVa/9AnRpAw9uTgDI6bi95fVbBrVMTkYGDJ
qtTq7yDXgRYL/3+St7ZUWVxJDKEBQs0J2TAl6qljalalBB8wWRUvCy6PW/fi33Phlg/DQw0Wah2j
0yfwr8BWw+KGnpQFywDEGEzAa3vZpKtIqec/Z/KN5SSE2xNIVtWBu3RQtzSCugEtj12/Hxi+8Tdz
BVHNGYtO7evWzRzCsTNSdbc3tWDUylPly3VjOk5deW37tlXOPkETbvGxEns7/tHQijgN2yiguAj5
6J7l7f7l1z7CTWGrIVeEYOiVA4Gn9lFtiagxHZqjsrGp4pM/YwuZaJKl3Ne92haTSNYZZfutc14j
lId+75k4NW0o0a6q0ISZNBnVJd2cqZqFKl94IAdcEMIMtIcmT7WjF6c3kjO2z3khntaJGe2h5uJ+
PHzoB+R3c8yVL+I7zFC8WNrs7dsq2qwGsQN8oVvatjSeW+VcCfYvGDTYACNXDKYXoHA7VHZ47NN+
FjRE9st+zO6ED3KR0+ZFdw3Mzi1pHMr5QmLS5JgU3ekCkepUt5ckpMbrUs9aMkDyrGRFyiH/GlZS
B19ckxWyMpFTl0Ua9TfNZJSaimJl0AnQKXibbBDhn7nKzsGnbnDBZEki2h73sWBv9IxdVi6mDCcR
tvfRRvXbj17Yzruyo7NfnXFFHjcavngi5SFoSPO5FIpD8YO4Jb7Fc+N2TDQguDTLBIEqyk77inn0
TO48/D8VvmUpU79QaKJKBnwbwtGbKvTS9lwqi42xKgqTQMIxsCI5WHZZ4VwsRTY+7KAKJC9ZMuNx
n99Ci7UZMI4MV0SNORkZugZMWyVPE7OSsemIZjEYe7oYsuoa3PZU8acKYrZGaVNngV1X/RBjgdJH
Nh0RNo+cJo0OfHpDy6DNhq67dpkQB57BaTQU7oNoZV/n3GUpA0LM0fs6uEc6giegV23H3FQ1+kTr
W+rZJ8YWsbfD0/GFeNORvpntEhrME6KsP1JNrsj4OZz7S+ObsqVS/kaCG9vIKOowSpNZPCdHtaqd
lorMpa4LS1mRFGHHLHoGZgQaxXQQ/8ALkaeQs+Hkh2o5fp5Ms32nJ9kCpE0fnxcaePK5biiXhKlD
fml1sPtINEXKukBQZoE5ikM8dYYAaYOM/OR7UzQC/iPUxNe5hj7zOsHfqK1pXZzvzj/OPxFY+8fm
ZGHNKQDZLgCarQIoK3fjYrtQz6Qio4MQHUtfb0whd9ORkx0KgOV/GA7b7rSG9XALGo68/U2ensWK
9Vv3781XJfr5clHpELuGlJMA0lX0MDBZ0S75QnLrL3E58ugl5yPYAOtE9Fdy8Djj3AbFETklecP9
FRCc3YVjgGV1veMP7vNhrkTlo8syoXq4ESUMGL8pCp8dNORsDL2g95u0hhCLdk1cR89J4/wEusea
MAAbMnttmYw8gIbA8kLs1Z+bdK8m2WFU1YTXx5UjiPPQSfqjiQJ441mkpnUmoeSVzPEbiTd+1iTy
RJ0CWtgnS8jtl+5S1Q1Ia5r87tX8Ds0BEs+qDuAnyCu3evnAXVZSkgvFRYHOvFJrMrqGVRIF1VRB
Q5w9Z+cKyjL98oN+Dkef5Ppbk9DhNFrDCR5heu1XXrX4lbKdV+5C5BsOzzcta6EHDVlLXv6LGMqb
4z3Uj+QsHULX/Cf+NmrK1R1NDqK7ffo33b9eDWf2cnCzT6MSilFUq0K2cNoOhCgwWKgLV430E6Ki
DU7O6mVwZoYVypPnp4meXzS9YulhbfctbYJnI4NjYmYDZ4CzkqGmrSsuOWCYuarkshRG/st9R8FX
iWXKiZXHnmW0+Ca3pZZBboE1eJop3V/GXzTCCS0H5UXP8RQSLtoFumZMUMkjws3cTcwfSzGMt9qv
SEsJPzBShiUO2gpmLcHPQb1thpL1rug/Vih3N6CsksA9xCMFJzf8Ajh4QqpHeU8KZAVcgMvSAyIc
BNLKuw23idt6Usbnz4EXNDPB2PF2YeFPL+/v1g8UajKp7+EYDkrRWeQWkWxWC76ZVZVFKRgIDX1T
KR8nNS7v9FMKjWqCHSTmLIrp3N1//nbwKOStqF0B6vGM1ZHB3KCmMn2v7OCDeC3tpvIwf1BVVK+i
ADvEqwPSyr4KalaKntj2GrTbbfsDXS/o6wbJcdVE4q1PVUUWMVRMYtlHfrqcoi4GAjuOQH61KF1L
uC2jt4yzSg3bbWGejW132pMWYzqPW4XdNCKXvkoBDlm8rvXwGk1B0jjlixBsT2SH60poJP6wC7q3
T4MrfIlLXP24z9YILL91OFmoS9C10V/vAxXpu9McZHc/PvkEuRxnb02+BD+vH1rA93trpWVVz7lh
adlqLZ2syv9FcvvvaAiAPbv1CiE1RJ0rweeJeaT/U0mgTU3Jpysmn/ZaQqmNUwy6lGjJ+yvq8H/i
fGvrc16kgeK9Rq1pZtJl97LBmHPl5SttN9wGWhRLoz/wYG+wSGCD8O7pd1x9OZE+zi6zYmkxeDFh
3+iL36l71jBeVA9jhUQMW/k34aY/h+YwuhS42nJ4bqVjbLHCbYtToyvVNKM32s5xH+it0jG8TLPz
AyD2pgcTtCv8JKcBwmva/gdKFBSfI2w6yHobXef3Hp/o7n5F/dRQ+f7waUfKEwz8sMDBzdw2hNn5
2Sl6/Y2jeWqG3rBo45HZ6nwFaHzuerW75pQ8auvJZ5P4xONf+PHKO0W90A6xDcr76j0BgmcWIQLS
no37pHvJi3HGC29+ynUayscpDHX2S7VkQHUIKtH9edA/ak6UFhztIiw6mVDD3d+gAakD6vzjV8vq
ZDn3AK117FGx3ZDKM//68wpKP0MrhTRV5vEf7odzJ3fuiWWTxzMXBPtDICV+WgX5pZ61vUsyYqgo
MBxwHMnIUWLGsq5Ch4bIIE8vRA8DSwqOlUqhH4L0K/baxDCm9J+iZvTI63oX8hFkFKfxh1zXA41T
1vA39E40tJodpYVgT8Tbq2klVkjobrliiUr0b2hHvxe/HZuvmTd2/hPtUxJK6SNeq8hwjkJtBhoS
ZTLYq3WyPfxkhCLoAWNQ9C48+91Chn1W//mboz/7mptHtg6IexWpN4L0xFd3tnUnbaiWQLdcsaMs
8whUm7TkAjZiwBczdQfz4B4Pa8XAXm3CYPuMM5Sl1UvkLc09Qca6O4p6iP8ac+g/6pSxwkqPawX/
LIGvQqIPenxG/fjiJxATHT1fYpZ6yBZQrOSX/y85M90ion6ACY05v1WeRrAquJarSSJ6Vr/TKRDI
9mVt8SzN4vtLeclnbtilJh9ja6Nq/j1IRMpebsBChRw3lewXOchP3dmB/3+5bNh/yMHIf5AjBEEn
SJwcSwrMnPwbTU1NnOzquU8lFjmVTwK1atxS3G38eFS7ypyFddj5RgQ0El2lzkJegNF3c3kGSTLB
4YdSC6ws16PWIh0oj7QPqOrE0qv5tWdITx7w8AvAlpZyChodXJjlq4kj23gPfrxF7sFk2R2nT8ns
OaAS2ye5PbRXLiAS8XoqNnV5BljDejHPppbIA7vJfXn1KruV8YWlzcmfLcCLtrTHZ0ykdZZLrQND
sA+to2Mfd38xIm/aJo2mZIAZmsA1kyntrjTBQBUCZyjIxMsILpii+zNf4XAkkHAMpGCkLm/AfXYl
KwEC7Qt8on2IH+cDSC7UtE1FKdOqJVghCeBOTbqamKgJf5swme0qj6eC9EtZqL02eFb2IMo33iJV
qUhcORcDcquGvU/sd2sQ0JZrj8HBmB3Hy99Y5n/gRp4ekHmlqWr2VcNa0NuaxDaWNKjkDgk4WVC6
g2WuR6EfRHsgdSkwNPkCSENoR+e5vYHgHoES8jZFsg/4YXnlo3NtZkJNkDb6g2mb55WoejYFh0hw
DFH0kXM6HRQ+X8EfGGLfIiEKcmr5qgHHdU/totAmUxUVb0FbIeHXP0nWLk+VnecM7OWIYWf9tHld
TdE4olri+LeY89A0g2GeYlgHw3YG/dMO+zREnrVBohoqULHY5M3kKSOkJYKJkocNE9qvmMBNVQi6
a4x4MhaWgCbip+wpLfKXLCKqMYqqFLqN+z4cfWOlDmNi4g9Zqx78yQa9tv+vxPMu9SmuN910ZYjr
QuOENFDwOLHWT6fVG4d246M4EUp63GH9ZPCucu8FLqODpDJLivcGJeJQqoShyxfczMW7qTjxEnGp
qn++KTwE+41t58XfqNB0tCKQfap1Mqca0+HTOGB1bwcGAL4obyVIN05lyxYrQ2DmOdb5al04PaTV
YvDL14I+ZfwKR2D5ZHLgvcPueKYRR6wvgsgNiPza+wZPYK9jebpaFFiwumzQ9G16xAYvkI5pJN7X
j54zjhPbojaX2Iaz1a9KyL2HLdiTPt47NB9+Ad4cSVomtRx8WrDqjG9K84ilFITJovIMqtPspapH
K1RmxvsVLLGIdMrJXfJ+PsK21GUnyAtgS+o+ey0HFRhVmd33vboWlhjC+Grv0EBrlqa4wBPmQ0sG
Qnt70kZTdwlUdM20X1kyTEDwmg60LgQ54j32aZW3c6E06M6HZG/eSblfC9Gfdem3xZgIIMFlwxvA
z3g2Emwc17cDPLJH0kuGOuJ0sm0kNHiG3WO5eB2DzFyvF9DMQnDsLsgpNeeJGr1fdpwDHHQZ0zE6
5rsA9x6YEgpW9+yRzr3Yn0WfIdjyb5nbbL1jjsUxg/7EdtNSd093w4IkupoJyo6IBaQrPuO1A0ji
fjvIjRliBlTS4NFqL9h0zCNPosGeDViudVULmsWrsbVHDaylQ2RQl9St227chAmHPLbNqZnhzReR
NjYEz0vM4pHBJET7UblsjpPhTnvfTfogr2Oy5B9j+zceY68ZEs8RA4RYtVy+0RJsxlPyPXSbE8Sc
t+boHdw1qOzSnZY6j6ZOw+SSuFcYGmHNfA6B72zuincCg8IJKLn3VlyTSo6/gvB9Nawg4fywj09b
9GD2p563cbEAhIMOq+/2qIU0JphHT/Wxk0UhsmQ7vaEzbbE+w1XslE2ws4QGjxPAzvi0wS8tvgS1
ICzAY/vtYHH8TURb/bAkgugLuEIO2T9OdLVvaINqX9gShk1t1dk8c0AIbSnwJ5n+WReTB/rZR9Vn
klkZhH4CTtjihxsWlollIOVBxE2FdzzkkMv8OEyHo/EyzG+rrTmmmTGOqKuShR7wAeI/TWGIsZnu
5JPlle1AuEOBpMsBGK0rI1dOyd8wT1vkvkp58wzV9HZwncEBfchbwy9Lm0k6xYBvZBvOOgm6op4o
aUQRxR7z3nUx4uVA3Gmsx0cFISmid71roGfOxHS/So3H9frnJyeAxril6BRG1yFEoJGroTldTWtp
4k422mLKIVHZ8PhEn5UZ3BuOEfR1CZWd6eX2M4s2daE3d/FMiINLYDkLT9eGyn+WTraOPvyR6tgQ
6BEHqcaq/jbzs//tqqB38GibhQjXUZbwo+Y+3qAruahoziAcSbDqRHqijL1fqyq2VRBAA5s0B6UV
OA+M9flItPvDrUKnpsAsVnPXgLCorXNEdy3ouGs9PDQV1DM195UARETzB2VdIwjmrSpgTGwewMP9
x2lt0J0Ica6Tx0YMU9JOVi497BcPcTH7CHKXUPb0LNGTcTp58r9jNDD44moGdQ7+NWM6HYj5EXFB
CMEnzF9WJWlLSR0mhJYXxXIrhZV/AU+Rb9ls7SyMHvBvcY576kPTURd8xUdxaXZGnfsi8cmrbIvh
0xa2U3oA8Ijtx7pf+V4lPbkU/Jstsyk/I+cZDbjMbLQnqyXYtrjVaKon2gOsPCcr00dOC/GWC745
EFAA/Aho4SOxklrsLZm2mDD5DxDIYVI3T1lhJE+ksP2VO50ebMSOFG2NCcUs4KxT4H5gfiP6FlmM
TrkS/FkubjzgUinpBHlswWgqeVg54f76Ouzw8MGMp+UivetdHaw034geD30tPg+2LN9rQBcfRv4p
wq1r9PngcUAebQGmXzLlBM8VKAL65y1DIpDCUiY7OLGcD83kMACt1rQfk7yhgjWY2KXibC5OEBeC
yytCEvkmcuFsBq2P4iPt0qJ0uNTanrluuBG4V56om4AlanzMHrRuG+LuVuVjOPYh9XhpP+NOHm+N
qisCFALGPD7vOj8fbbFT8Rn3fXtifVHc45XdoiznUETLVXySAI70/iJRylESWDsorhK8oQ3uf0tk
pL3dOoBq13Xm6RttYxgKnkUzre+Gn+PBjepKRjymVg96RFeDsQqnfftmOEIJYozBeCHMITVKw/AY
55C/RHXBihWGPuHYnOviapG0VXF8gJjM9OesH0ZhmvTWfgCi6l2wzEk8fzkU9tuSsVwAHxsYBo4m
b3kZpTER4oKuZynIRKts5X7kVMkNT09fpb7XdLxzIUeBowM4LussNWMlDIFgjDnENe6VEhcmxIBm
BPCuY5IyTzaF4rBTkHSdMIhkr7FjIWaZIagqOL1O0P5jJ+z6xK6uEY1HFxRq95QQCJOMAxoUYphx
HVqt1RGJV7kiMcXENkxDcL0/t7k9coPTWyslvGHM2jG0+DRFh0469vdKnf8QagFY9xFwdxLtgJ0O
OJPHN+iEYa78O9fyQygVEhxilyvZhhMlEpsleL42sJV1pHil52uiegN2QpMBWJzIngUYBCAMvQ3R
u/gacdqSGPc109bwWSs8fHL4L9wTBFMOicVNI9AdhC5hoSzdYJHON0XGzyvColhJ8IwE3TDzdjk+
+Jqj9wQpCUMX0DESsJsfqeqdm7KQby9lVCxTMdbVTICdGg5omZh1A8OwM+T4caS+AdCvyc/k7IjK
SQBE7FHrSqXpd4tM1wmtKdZ7Qa9D/9cKckdTh8/isKxY5dqBFjt7Y+iiCdocSDfAH/NmilupXZCx
UwKiEtVLiN6NensN0L987rLLlGK9OkcBbJYBT4ajFH3Tbt2QHQdFq1vxBK9VdVNCMjN2/axx18li
v+lzdstmE4k9zwcUhIpL3yRxwY7ZbNdAMacBqCttwzJ41bRZxq1Q0m6Fy7mt5tsl15B6SZlUFNtF
I7NW0I3NB6IPLz5Rl1Uz0XL60io2BE3MwhhB0DvdNlXDgP7TkTfKqBckmK6Tfiexi737Gty9mkkS
eDPr3bUTcDeY1sTWZ/X623egCYus7JAIc1aP4vCYM3FMBk/7wwYaoXhrMNAFUr5CJ8pp4uI1CAPQ
R6FRewOST3RUe+MCjCHkiMWBKwiMzwWWUOg2/CZqGlHmVQTo2hLNxaVpz3LF7Fm16u/PQ8ABMNxf
yTOtzJFYef7jt/qhRI7Sm2I6S/vIHju+pfHTDzGrjJQVilJXctb7/ujODhQgcJKRuG/GCz0iWThT
05VmpdcLUHYxN8BP3c0aV5oKUBlpgnxNboeVdRsXXf2vCYvi2eHzbSlXs9Zue79wKHgyihBWQBj1
dJxiMYhfBc/1Q/zs/7SNGN7qjHz/SmdnFrEbk65q7n+0pVUKqlKanxAtHSzyZGR/iB/XtZWxKA8k
MebCQeloA1LtF0bwjDK2dUzdcrWQBYBhG0AsUhlwBSPVeQHtdt7pR0oVNYucQXrOvp7dCTmi+xKb
JGn5Uri6ZvRrBUQcQFg8+uic8nRNiSEu69I5Tjrxjl6EWqCK+AibcXXd878vkux+FyCLnvDBINhB
NrTpIwx1+kB0McTkIdCZhEPpogAcM0nsfrdQeB+72Lt9U+1AlvbDIm28cqJhGleQihE3R6V7eiqc
5+LFKbX58TBUVBtfUCM8gg2g6PZnzcCa7PxAMVu3RbHm1PJJW/bsMvL4id6wsm6qe+OUo5QGVfXZ
mb7I+Sml6CXinDmRDoRq9dw5+BUueaHrrINtQQPvN4WamrozX4I4EWFOcZe5BKBo6RaiL/esUc1L
3k4blu4hRCedbDLdhUXBvq6QmpFFzeZn9WQUCNOOCxMA8Z8NvlMaty6Oj0xR8GCiD2pVHy9POxEG
UDL45V92Wjd7LxwOgAKajzO6bCg+0p2eunZd2D2LbcGZdSM9wm8fove/PSMJ9A1+D2PioHJFoTnA
5rzF5UFaxkQqhPcxfNLKVzMVW9NrtdKNeOIP+bYzXpAmwQC5/xovidtbArI7qBivSUEUaY9yw37R
jYGkkuula8kHDBsrVSarQhe7AKd0E/LWa7lDcMCO3sVAQM5dmYXhQCewuhFD1wqvwvei5J3VKaNn
LxwHHWBlZGOyn+Zironf2O0rRpD39xzJknMxdm6aTDINRs+qNtA3cfy0BLlabBOWnyWjdcY1Ix1D
3V+PlsHMX1UOLfEztl7XlpSSeyyfw5NkfY6DEYjM10LEjAA7RyWfnDeWwWPvcgYU5ev8NL6RGa3e
pegTzN9tenHEz8LpWI5t0sulerOgD69BJoNE1UfY1L6hssk7Mii197Iz65QOS9J8jwASOXdf0iV+
ixpHIK5fFYPNcZwkD53/oW14vfkk5rgzENUrFul2ChikCt2qPi1v5PD8I9AEyrBRTVatG8NjlwkG
Bt/UxNUjpzh4iQWtMWS7gnoCyPpspVKAWDMI6XnDaNf7cM71DXlIw+PZlLTLU9mqzD2RedbHY26T
TWxEMBl4xZbhlx5ink/kQMoyuG7mCWiFJpPIn3EFTc4XlprIeXb9Icw7An0cmUkKbxfVYMGJ7ycH
qQR41E/iRTdHDiHV3VTHPpBp/v3d2F31IeX6GR+KRk3owJFoxS48nCW3cU35uMr8EDgB4/al3puM
yTvu6ZbRhmdyc/DTeK4TBZlZDtQz3yVv4A5MPQOMiv8EI52aQBFT46FyeEol1xMTZQCLfUZG2WXV
8aFSTajIKGNcEhAmWRsR9mP9YRhgx0UMRsXYolj4Nx8l0MxXK/uuKWdflk9Xz4MGY9e6ufPa4hiB
kWuKqaJYE8hSIzBZ35FZ4ct72Yqa1oPIC8e6nu5ugZfGmmi5cX41AGhGoSzABLcdPDGfFQmYJYyq
YrXD4reZfPGb+X3OJF5rM+wQee6QCwrI8zV9/n6oJeSR7tOffDhDx7O9OpN+kTgvV9GhErw6S/WD
LpC7LbthUl3EjUx5GZVz0Krzj6cS/XVEqMEfUsZ5W+Bon993K9QGgHGvtTdr6fw7rghhATqll89g
WjUos/t4Ug+YEfOyz/NHHj1sOzvWIUlrkqf9MoNOUJzzUnTaHvEf+eOH8TrlhOQNQJeTb/1jFdQu
TnuXtLwO8n+ONbOYcPGWQpYQIZDK274pL0XwJfwQ0KQc/O/9j5fYiKwZ4rQOpbX0x23ROEwk4Wwj
EO8aaG5mgTBrhu7uNVEtVEfZVZSjK9XnViQp42n1VuMS5B6jyyk9ihnlsUP4rl4p1TCIxYPhTO9/
Wh7goZN8mRY8HR5uBAOoNgX38p3SUJ/1UXULzKZ5pLI7CbZZGTMS2MwO0AWgPyCNiUThwmVYZVBt
TrlGe36Wf9/VDZJ3C4XYjpgyi3AqANiBiQWHAu97E2vtXj3IwU78cb93XnvpMm/e84iFGb97G6tT
36Hc/MAfVao36GCDaWQDxo/urN8HDDGPuYUgA6HkB7xU56Z8hkZLDKmmc4Y5rDD1pUE4ZB0NSH+Q
PB2R+MLBEImLjkT7bGoUdF5xDfRnOxl0DMIQU5Zpa6jq/1PQ/qlcCbXb2ANpwH9OmkdvzM3ZuBdL
eLGi1NEqCD4Rf9gEYqXirMcNMbT/iL+Y1XAEI401+7ump3axJ8kJjybpmqEFmJMvA1Ldo91jc2S5
sjcigx9YyKZkGRVKPK7UomxaCe5B1+j6jg6DCPBG7xU3PiSRuv+qzru4DFc0rVbdlHPPs6srPmpu
CwWCLa4KMyuVb5Llgpr8MPA56Y/YuHzRh92rIIkbDQw+vh+ChpC+xW8+iUMGmQsFBZvMvCrOtD19
UJr6GWNWWgTl9D0n5YEmeF6QQv0dqeKSVRBUo5IxCR7mYNmBnUo5j3oNNt/Bx0b89Ooh1JoCRF+L
d7EtPts3Vxqo5J14/aXSIQEgsCYlgb5JxLs8ZOr375jfR7T+gK+6txYSxHxpKzHv7HJrYpDpOSgM
vlZMQlpjkyPG2pMmQPZBrcMbAaDuYZSBLCS5cxAvsHxRcLTSc2VgYwP3YDoxfHwKYOW2VkMuppjC
EN1fxMcCUhDijCo0iY1Uy5f13wBzCBVFyXe04lla4Vg6XPkpMPcwBTzrn06Jmi8H27AxmjFWn6iq
Z77cvFXQYAm/V9ea4Kfb8EqbrOK9WnbxcDoT/FueUccbpw3bO0sICwnTtFMBxoMzKtR8PZea/nOl
HRZ0BzHwIGm5YntMy/Na8KmIJufUrTV30aiGmVuOXcRPIMlf6TiOb9tRO6atFT51VlsV3QeY27kp
NyfAfI+wsuorAvIqLjNf80tFDRMZIU4D7/DyDZPdx3oHTupbbXFr8Le1KezIef29m8A273Er1ej/
qJPmJY3BAuDtbYYXGuq8KkVhzScl3UJy+QAzLGSCDWhQjxcny3DjA09RFP9svPZDqI7p9nXlUI9u
YSIRDCEXbR5JcdNl4TVAk6zWdvLW/8qxNc9/KIOycMwY8ZrM4+8286hiUGOs5UgV40cGN6VKLWVK
u2MdXB8mcIdsssC9ZYFU1aa4OibP4NBEkQ/q8x4A/V1OjGIF65vtH2SyIQpS8rQNOxaAE0YngWi2
CLD+0ad5UVRvxwMHMI92ET+lrOZWGPk1KtUanVwEM2OUq++rp3flkrLnVY6654avU9Yk8IZrG7oK
0e3fUphhW8DbQmbCbcC5Ib/p//v0zK4WnaUzP07Hb7sG6wSN9AXN4ZeyqLuYA2fRXj4fRURnnkmF
6Nh4DDcCg3fzrkIeYYNHDuX5LlhihRT2t+RlQ6wxtRvUl0bZ3BsTxzsefT82XhZTPwPSL0v9Lfa/
ub5kTNIv2uwI+xAbtJTW3teoksLM5jGgOjKFtffBMGas1eRUll9ufpEpmqOE4JpvjmTuyx3wPByp
W7yBb85+kO7YF33pQwZKkEDvZesxWq3R/p0YtIrqIDV6ZtAtgaHqMnDQvybYoyo9cq1CSsvaXCYz
sJK9vXIzHCnKe0I/WouU+7LYshQpEHiC/uiFLtFCsUBGvkFyT9IZPU5swapp/+p2s3ySKYv5kps2
PxCuwRxnsvpqMpacUU4JvrUs937ynl/gWLpF1p54SoeB3y/O6IhKJyNM38lgdB7HTkOma78Q0rzX
Wsb56Nuvm8Gu8EEeXci8M970+eA43+4Mkd793DP6P8vdFg/dglMl1QDlUjYlfu3iZ1mpwIeKdaPl
v7I6QzdcL1A66MFxIOn7KwtMlmoYs0wEWyaQIPfiAPub/4mlsOh4/nzUo7puZhMaOPyUcMZYLZeT
8kCMvgsmedgpyVcZYnfkOidNNMNOTlKOUm6C868SxISxljdG7g1Baf1z0uCX7+QbxiLwmUwW5mre
3GgVNfGipSszR8p+eaJVOY9wkULz7TKP+kQlQAONLLfz20T/8v/8+5kDfarTqFOb7mg4+Hd5A1RF
FO/LorVhEZ9VPvc9dJKDbqs04Zlx7VDGkS9uYOw8d+boqenho6ucaAxguB1XrG17ljw/g5er4nmv
nn+lHuKziLky6YmGpev2maOCXYHJ4uwRi+v2PepIz4czmFu3LDuh/PMRtEwY5aRjrEymD8+/p3b7
mTyQqzkPfcTvMGQJ5yfz1dv6/d2pjqNez9UrGH+txFUIKyVOiNP12Ik/ttkqrKX3oq2tR7B3/THs
x0UpTfIebTnicg8DzDIH3vee6qAOmJjPJsBgxfnHKMAyDsLUUB6iLc1NT6JMtjrZKcYK6EV5Qdox
EMbmfETnXMbUUdpFzRK7DZYZ4r/2nxVCmYZnt+B2U6cUW+2IijVoiQGN5S9CeqTneaJyW1MaMRQe
9VsgOP5Fkfq5P9Q0l+28Usx8+E535k9LHk1ir8k/vXLWimw0aCTuMw1z+LBuMBVk8ibMK0tMi2wK
uLr/UrY9j7Cvcu84tW7yq2XL8lXKXjFlHiUfYLu19NOoNcwK7gG7SZBZelxO60V9TLCo4XdSHPOl
fkY0+pH5r5mycwx6vDgVpFDifrKGYz/E6aSxbLlKs93W5lp6vBiqwcEONubdbnaRdK+Hys2uZ/zg
XpP7fDPmU38nIU1ln6TBdKS9oJ/gxGU6EiPL9rco/P3zw8DwwnCf3DDzppG008YLtRXbyK/GLZgy
NABlXzm6DPhhUgZgTM8Uamf+5HpEIzza1OofHVGj/nmmyddrSKbnYKasDE/89YOzmX+soL6QTcqe
SCY7ePrvmCpHu3MIdGWv2sT10ik/0X2m+SMnPZbk4t4ovwPR3r+EYitbMEDPFAmXjFefHWt4I424
7BYv2fGzJ7Bn3zKWbgc+wsUS5D1JqYRutQK9yyCFyLRgBd9dl60BrwlVy0Sf3YSa8LZ3gESQb2QW
Y7SoGpjFrobjosaSBXyil6YxVLkL7JfA/0KT4xMOF242DGSEmzdm1OYtQUZXMaZYcv/O0JJfvgbm
6yx4tZ3VNT4FoVnH/QKxEmeSu1LhBNtK18i10glGin/E0svUTOIXA2mWlFcirZS7IEaZOsep3D1n
W0sXR4MmZechf5w4rQgGXm/WfjdkCrsba2wx0I21/VOKbrQ/O9BZ+SpJcVCed/TN/bh5Hr8IZb03
s9MPfTqgue5qxdbFMGqrW+FLlV/l4JQlfwDxO079CyA8M0/kfb923YnJ1lEUTlrml52RrdCdU7sT
xvHaNuX4WRuyjZFG1zz86s4z1WXxBpLYscJcHj+zCpzb1GbQposqGGHo8yZERsbh7bw6yXZHNtHa
JYWELrxhvHifu48AIZvzWNp/UCwKsfVArJWmedls8xsDC2oU5z5tpUJDMiYrF+GwZdrscG1lfhNV
7kgXJgkbdU4/QNTx5jLsIqeW0anYV+P//6wWive3BaF04PsEY7x7kRScbhJxZPHGvNyvHWdvlhUk
pZK1ie+k1QP8tgyJVnHdFI0eqStGCpo93jsidZxK12yZTVLgvjUeaAA4jLkVse+lQvGkUN+oyyt8
koq0zpomtbH1pvjixYV8ahb8OPVqX9aSUT+pCpoDvet+TMqXL10lZHb6ek3S8Dhlh6h9NDFELrWU
HxlKQCdxxZhP5EYmzkQVYc0SqmGZb5gEzAiwWaUS8zEw9WlGobl56OAaDtYKOgOdiYEbtEYycEa1
+16xYGdDDAu64ACro8dtJeaUWEhLR4o1u8L4X0eVyHZuQ/44LEm4Sz2DqIxqX6JfviiAw42REe/8
pzJy34ERXKOUpKY8HY10TRVQ3yvXhon1skWodT94uS09XJTAOTN0VhLrlGZLCk2jfx2VTE3uATTp
qq04DbT+TEjx2+8/f1FtRqPaLvm7CSx3e6gn1jEAA5E6b1gNltqcORu25uH+UPSE4DNu+84pRIqJ
T1TWASQ/YO+nt2AW38uqEJy5390XBwCS/vmKpcQ8Li1kjOTA880WxHG4IezyBGyw7E5Fp2j4/fjn
4/OsQryv+ti2H63ULuXGJtp8XJbDMm20FvZ6ojQegG30fgDIHlcdxcCIO4Av9nP44pUbNGdxEVC1
EeetZ/jd9Pay1QAfLlgooVJ7fDWaTbet6XI+q5wgO7QCTcjy710F8kz41jjgmz/2o3D5j1QdN+Dn
A+bXyToSyYZfAJvBe6RnWbtDbw+RTNz/JrklxoEl3h9/XpVqdGPgN6f0PvaJ8aARpPPHzN7nJpGU
dgZsjAbR37N5WG90knTGXtLvKut447N3T02YJaH796DxfwE/5YwIPlLigYeDzDWxwySOXoea+ESR
O7igR+l6YyJutyVvsbFsRqigUXv6cHaWxefZ9qDffeqyFtpJv0ObK56DWLGgfcsWkCdife0bOFh9
WuwvatBkSXTrr5F72XPXRNsMhaVAn/c0VYBEC3tdgx338urLDI/7GpEqVnqiECYWYU0lrHT8k9zw
6KQp1zn9FhMlE6cSKczm9hop4mbvrrgi3XbRXwlQpKxDAanoMr2j+UAobth2IWT3vGFLdE8A8clU
8h0ouzGc+MMgzI48i20SifjEH8BLruPUHbO0Fs7tIyX0WCzb6/4/QV0kf//H/HwU7EXk40mAFlC+
hEbO0jeisgwkE39DTEWn54TJhJCZe8BqPlMn3l/qr78VhUFKkvf0DpAX/bnWnhuaOCxXFsOZbjrB
T0yEVR8hXG8pGj1iejMJApxTuPMuYCpsIIunDjzouXm7YNMg8nEC2m8wSMOR+3Xdk5Gy3aZbn9/A
crWdJ/rKzr/1LG6TMRZjTWCm+coLt9JWoo036KqHK5xkhq86tnKnsKRnjCO/Uau/1nCg/HmEfsh7
nWjQzu4oMuxfyZ+Zc7pnwo7Jr7iIF1Zh840ESOc5hYjXJujSG4cb4nzfi5Uu6fnH6D6QNFXFcJXz
+NN7XFUw6BxmQCQk4l7kTQMNYOht+2syJMCVIdN2keWK0EBirGyUv/vO76F2QvWJY/qfQxhBQQvj
E0RgtP0sD9bcLQjxHSK/kCuK1XyTyfgFw7wI8Ho83Isy/raFbMXR0Ld81d4mIAmF7bfIqAlsAj3Y
z4RSNQvI3ZgWuA68A7sgcpl9b2aA/qVlcD1n1p7DHPbXcQllLRSnJLN9kpWs6/aA8DRvdkJ3cxGF
P7/f6TH63w2Rkk6SC7JFi1XL+w3tSwRt8qHhLDji0C52Vc0SPRvOh7WF9Ng0U7amMS7N7Ur/TD+T
BmOLg1GFqz/erq6eAF7tKlJVENtGoxEZfoIJhTB/XDjghONIbtqgxXoeThOmg4RttUIl447EHbbT
Z+nUYo37pZssim4PxiiI5PNqrlZf/uJithWBpJLmg+fxTpJPOamam7+cxaH3h9Eg78guzJfhnjfr
7rMpN4yPdSThUNAOyFMHN/AragQ4MXYR2/9MHMjUPUF8PuAP4VfzJ2JQcR+fevF/V7L13vaP+f0R
0xeE6VQmTOMM/yaTCT78Iry4cdgH0LPM3ymYyHM5mHwbqM173mgBVqNLCHFLyPSDIEm3/tEZ7ocG
bAnuFcreSxL6dNdH3IomfooUvqF9zYs5tG81xsjfRP5+bioYmRAGARxy77IUGBiX6oRlr3wEf8nf
NoLpDYyl8WFkxQZFCT7mdiAs6IlU8y18Ozk8wZiviWxJOfuRP9fvS042TDcgNdP919nJtJsKaZ3/
Uv0cP7ffCNK9e3loQyn+cMGtF7hya5h/ofn7ESPZNQqBkQGfvmT51tVebeU2eZ7+zgKKjV5Lm6i5
SpE8/mCCtMrg9S+wQpaE1zXP5fKhChSfWVMNgoQ4L1MIrBvD8vQh50aOjcbfk1NDMDhODsadrAn9
/ZuAs8eyPntV6qv/wME9ICJ0lw1Dqob+ht7XOhljRcAMt+VMoueXLAH6MvRA1NIULTuA4MjrnaIW
fRwORpNkCqFc7jvveJX23IISII/47dZMTFjp1XDK1l/5LjSrggfkyW81oCcsT18dNflosERKr+HU
lYo+oBoKijj10jXBStfI3z324DWcAKlWRcoI4RqE1qMei2V6EI7q168fQHqBwm0o7lNrkLRN/nms
qdjuBHG8yJMSXlLTRTQ/H1xSmAFIb/SdBNSW4GRSuxQGA4c+b3nYiL6a/42YFcrLbRkMl+ZKpeMF
7g8WvjqcATVftN36/OeF+KwXtL1ChqChznAcdw5k6IXij9rWQCrQ1ycPSIeNFn10AHOVI+wfrXlB
UHNo1y1JjMx2Bp72KwNkrH6Msqw8MyEETVvwyXq4cEh4V3sQ/XZb62LsvxNmL3YTKC6qu2cZ52Pm
PWTy2YnNS+2UHmsMM8+V/bO7FInkjWT7LgHCrx1QJbWILrzyX5ezs9+7b3rs4ZKfiRAtQrF//zJh
sBQW7TTzxRJXOq0dAqji6dTfZjBS3nj5CoOZr2kQSQtfNrc/PnGgey37KkI8C3WHVfpC/DZG93cW
CnnhHTHx1Uk8l60bTeSrMjgnX8hVD1hobyh7LwGBj2Ojqrj2JG1NbyW0q1n4N5ZzwU1vyQOFEprN
SGLXKSEm8eZyyfoxzpYhVYXwdLzGLGrp2UAXizinTjACjGPs7llzYvGQpp+Fd1CAp9vfLqsbWi/a
gJZF/Xr0YEohz3hqW8+aiLhZiOynon/6L2tkAPebDi2fs8SwySa0aCL9BRSuzrRobkcHeqUBcD7L
8YmQgpYNV+k9H6U0rUr5oRa+UNTGtykfeQsanZ5xWgvjEvEpW6GSWGty+cFA0Q+/Ua5r/7K013nU
d3equJXt+50Bbguyxy3MbhTJFtkVGI7PukNKS0jSBTLIEKXBpnaWwwX18UPQ/x01oZSHWoM/GwuZ
UoV65LprzMuL/esGrxt4ja9FDo0w5yKfuFZHmb4NE62zHsKT2UYBaQZB7Ua+BnRsKcFa8kQbRVgT
trWzgoSKDJx8Z7KHTF+gM2caEFjpNY4DsgJsvc7MrL7w32zVyKHXbwc6xM7vy35NKNwMH1F53q/E
bm7G6of+ZnHha8KVd+HRG3vQycu0OcLRBE6laS5NfmxlhC8zzqYsWWQWbV4+/wiP1CruSuOuxg8t
KS+0fJEeTZBBfaa2nyEqXQ5NUpSCVFy84Po3fb/I9sUc0Mbcq57wjXlP+mdwfGjFRjfFTqSXfHfU
idMF8/aa1wiI4sa3SnOC5Id1pI/3hNaxAwWDtv2oUHISzDFosldJ/z0N43P6+IiNDzSodocqGRrT
cDlopoJEEUPcI/+m4xNqERXtgPyFEkHdoDdT/5Tcur82AYNvtoTdQo13ItRheHMNQmUXk9shcC/N
yY6dd0715WZDSX1mmGU/cnZxb1tXSiq7E3CaiPoRIV9sM5rLNazqXeGiu9v7UgVR0AwU/TK4VMBW
VHNw3EcJDjoa7B8k1fhQCo545xXT9V49wSpIZJWp5LB15ewX+yQ5X+JmXztxdUT7a0DlCWxeOsmB
Tt3K0lT+GGwHFzWfeuDvH8TH1nGGbxkwFdWPX5yNDQxX+o+H7ecJiKzyWA7U5TW2jGuvxeN3RSzP
iMkSDFjgLs+EOvEITcUrITcja2m2Q1vnG5CQs7P+Md2//h2KS51DdYkLKkiMlJB2zIDnQq+tB0js
fQ/7EuES/asd9R21rrj4YgjwUakG1czmVOk9ziEq7HQMahX8AV7c+J5f6tdy0nO5ACkAqtmGWJ4f
i0RQVJFXLKQu02rXM28QFUtUILNuMaGrHiEmeYKn6ebBGWHOi5+wHm7uDOP6suYJhrZ17pqiF5+7
pXQ8+KDubpTl0cMplqSdei5WeaMtmMJd+p1xMfb4sKjmKq4ynyEehPHDfzKpymKis2jzIG9N15jN
mQRUCQxpcg0PKVzu/pSMvsjJnA4p+ZoTeuuW4u9BF0DEaT+/14jHJmZvv42cnHcQdNEyI4LQl9Q/
zXcVaDv8FM1pciSDuuN7d4pIJhrsPcEhgaFls5jjMMN/6ghYEjO6BjgpwCpgopiTwW4qhCkt096s
TxDFUTuPLozv+McugvixA+okfzKIdPtPcByvE8iIpttiogtjtgO5pBZ4FPFcZWqSiup+FVDviGpa
8C70wmcp6QU65ywgG5uXjrLI7qDlf1kSkgeIbzavlkiB1dqzI6w9xsip7sRdwbPUTkxugNhGwC+G
9Z4XeerCYnBtQwzTHVXMyu1EZw1MJ1t1G0aN/oNXHVHUpZiJgzkKMdijMnJRGdwazi0B8Nd7JUrC
1aJw77GeJZxwNx+JJfRCatOZli10AYHLJvf+aLv5xTLLyJ/Gl8edcDM/8SkbQgozmcSccuSgjCF0
C8+aPWn22sAZCpkDRP1knqtDL+p1LHmXuRWFB6i4rSGDC5stybymM18l1fbF6Cn/6kYS1KOFgexZ
Nc07fh3o7NJT3naqm8tiOaQg09Su5MDH8PsxJGFDUIc1Qw+yOMpvoCcKjqNgfDud3bwitm21AWCB
iOq2AOMZaM/jJoItLVbXPD2f0Y+v4o8JICJX4Vj/QZsh18/xWM05Oyq7a9+a80gshVniC9Nv6A8j
NY5wUEDVSn063DlznIplg949MUGJCAv1nIN0OxGZZvCqeEtRvbrzse7Jr/+7lAUdFAuSd1lDSl8r
huOYYRsBIMH9osNLvS53lvL0dafxvWlz74iBrU4KFIehu+hGeub5quUsplWRQSGjTEIRQqsiPepQ
K0rmBH42GCckyAzsZnemPu/acBACLaXTuIy/AAdeyHazkFtdO3XW0YQP2PmlsiDgdSzseTm0j4JS
w0u5hNj+E6x6yvFNyN3OusMWHoNzCE116v4dYRt5kCRcmrVHHDyKLr/+GHaNg2LHLc4fUsgiNUG+
o2O3eYEFC0FRR5B/LrQ+INacsJNvnkQKP8YlhPx7wTOLcNd2AMrrnK0mELJkPqEFKCkTN/nnCNZJ
etE3DpH5tXG3+MMJOunQPqR70S+qvqAJqdJtfNG6MCWigJMWTlG69qCG9PBxRO+7/iTvAShMe2+t
c76na6BEdtu5VScsh2HQFNB1p0xlc43sY3vyQT8vb2U0TcadvPBomYN1L58lg5uO+jsThP8ZcSRg
szBK+mDXlvu0CodAbsh2po7uSjLiYWFBytApAGTn6nKAIRXoPPE8QC7ntZnO+JoL5YdOr196Y0rQ
xwZIb3QvhD6lkk43YEJkXedvU1IL1HPIuaKNIVWsTDTX62VsYNAuVV0rlWBth8vJBZQ90TV/apuR
t6ZblhWFCIWa9uYSBs1f9IqCP9raO/BBipxSrCRoQ4smWrz26QL84XbGd+DcLLvneRuBeQdMQNAK
NAYnW6odcQdP367xlcw/CHFHzWC5ES71pNGiGIH6m5a5o2OTBJqMw91hp3pKbNRTnYhvrFRYW2vL
GUzyQYqurlkZ32DfLoCflln1c9UFS9eCOdpuKLSjN+xyAmrzs1OvGPClMga2D4LiRNmzabVEuzZ8
7MuPeIEmjfUi3abXg+Fa+NhFhJBfopG/qoW9SUAgzzrA7k2iuGfNWCbGqnYnkHZDprX9EJMYwSrm
TRRCC+GiFYbuUwd3//vcP4uRTGgKqNL/FpgjSXG1syb5H8F/gH0FqIfRd5d0wKFqjT9ImeR6KGRT
dHnP8OzLTOihD+vG22xnAZZExn75Ha+tKZ2y8m7Nis2BaO1B6pPdJygUUTYO+gjfmWjFh9OWUhKE
YA5m9O0eg5Bfey8qYaR05+jgozx4v1CW60ebAYcr26FYWcBcHmOJiuAMpMXZgCux5KENgWP08L9F
PtqAW4bmX0nZYHUU6yIHPma6TtkhrPbV0LGMiCzQv8irFRG1/u7VavJw+/7i2YBYperBO/WXO9uq
8m1RhqKwfgQR0pg8xr9RkSNMbsL6etfHVgoso9cdnxPkNm+D8naN6Wu4G78dcQyL5ZkspZWpWl7H
YwIvH1Fwk4FYUn5Sd8Xqvjyyu0UmBre/wSCMMHaheqrNlHQaRycWN74qw5PY+Tl3zPSCbI4Gv8Gn
Ya7H3THj6d7xNMgZUOr1SiXkm7jwIzdtv+j1h3knqfiTkgeFqTC0KFLRxK4IUI96n1k9RPQ+w4ME
hpYV3FztAIWLBWFHdDxDz6xRjds5DYxgy8UqmZLo7Oxf5ESYKbQbKK4bs+lODcH1mL24nmnPh126
hzItjzGv95B2VJtuLbIFH9KeUUmcJDaRNnaB86xjoPg+DwedWclSnJvosUbAPvYtt5DLoCWNkv15
OvoV/aWgn4ZukBeaneqoAWGZNDGZlkdQptLV+vWzCoAYgb7sA0KK5eUfXpEyXj42EONXHSPmQfCf
alPgM53dZsbI+stiHfUaa4nzrXUj9OmaeB0/s+oJl6LrbwBdRPzZx52RYQxbLamH1r+fzdggNPjN
/VbYDKO8EvIjYvaQj7bQ/jBD44egsourXryEQQyvp6t3T+MO1JcoEUhiQWtfds9QB2Ciz39SlkGI
pkCsZYP9I5dInOkXt2kjQ051buZhQbPNASHPACo6sRhidu5hPYJHSNfSYCqsZUdtBa7OPPTf+SYf
w2N6UvuQJcGFL+AEd8HvJMNyKgeud/6wUuscmbrgygsnZxW9Gd3usOMHHIwHPLVnGt4IbrramuBL
ldrcW3J/GSRDbWSd9zYn7PRDjOpLL08SaJmnFbHoNOZTMmRwkn9aV9BgW04wyt440Ath7rHGtYaF
s9w+IjroARi8mhE8ytfEwSbNkYXrXbsOjK4dOTFNZsVfvW89nG8NyLOAkPvGEekEEDQ1Rs9ofukO
Fav6sBTmpnF24APPuchtM6zQCm1JNEhNtR1qlMaGKlt76wwAnme7+FZMke66EIUteEZeISmb+doC
49u3tRzCvTHR9LWiLpL8/htXbuui9T8tByPWQnbPKLePLUPYll9VRRqPgZcv+lhiaAuWq8hfFcsV
gT42F9Csf4Lv+KbbdimNxWEURCCUugFNYEbwcxHRvXrFaJgvX5XCnL9yxWMlj8gh6pzMnkXcqov1
8CtfIB/QLbmdmnSok5h9oHzhkxF5qg6JUffy38Hl9D+QN3sonOPK5jXYzUMlmdmMWGJfKXHH8Y0j
4n6kqv4EWsD3FGOfR3qpJZor+bAYGm+cYJGrc6byXrGHhU3Rai7iuRfrMhiQOZStdncMH66VIEM0
0R0opkuq5S8Hc1GsQDbuJIaAAZQPSfi0IwPRI3sRToT0ojmSlGcRVo8mIlpN3JPfHrIokYML40p1
GRZuXPb6rBt0rw5DMdj1pbw7Fy/WKBpz3k2t0PjjmKoJbWkzqzbJJaf3CtvkZUokf8p/6Vaqrbpl
yDX/kNEcLDfydkigbBQQfpR+XGqFfvVDRpQRaRbF+jOwlK61mIZODoE7Dc3X3ndjOfLKJWkZTwWK
SmpEw7wcIy7gN/8aE2pH39Ye5XeElojxdtY4ga3a3YqNmxnxxX5HC2057tujcCcU5d2eC7a54pSC
UTqDdygH8gFSvTjjrhzmdBFPCBwEBlSovrK3pwNiPLsHgIQF8YsHoCgoxCYYEXraHGW2fb+LMnq8
AzzV23Zf/y2YzWD8Z6qFV8IVAQ/CJS2Ys7gaRhR9kN55tKe5n5K/uGLQIYgVy974+mAAYBOPg3/G
lLk2Q5pBYptTKwAj/a74rFQnMVhLNmgT3l4J3Be39yNxiBhmWxgqPLizjekG6i1AWXP21XtIWtU5
HlR6r4Sf/VFVWKF0dSKcfxrxWty4uUHvI4+2fjGpOdzxQa5kZnJH8q9uMDeO9L3FEkJYzg5WGE66
ej/nLBNrgKKiqCur6TDqR4RT5F+Njc9zS0+i/nuByE7Cy88yShJTi7sBYCd0lw7MLpeHeAYOkMTs
cnrVQQwfQWQ33/KZGU80gkUQNcETZqRSJqvbwI72k/SNVzZI/tuqV2r/NReG1Cm25MjYw/XdNCZm
JqT5ohH5j1MEnIb+lw5XedRjpLc3XTjyhnxWm/4olQR1NnGBBrTyrfZ+lnIjXW4Cqh7Znq2sjc8D
YTO6Maezjv0VgvmLs9paJIQmOAdlizJcy/h3a4WI6OmYS5WnUcDnxEnC+qISEtFgO3UTFh4xRCV1
GSeinT5hpc8dCA3iJAM7VMAIv2s9wLNLqPPptQdur97HKm6uCZseZNJRMSNNlhp9yMetZE5IHBt1
dfBMxZAzJxFIt/n/kD7rI90rLqcPK0ATY6ZV36s0s6wtyejCN0f2SLysFSBUyXq12ROq8QMKdEqJ
7sb0cnbr2ZgM3iFndKrRfHoNTOhIuc4waQ/FXkehQlqOiiXGT2UKVNA2NhKscjLWrdr0kk7xq9Cp
tilw9+xlDXtHMoK9EJdZ2yu7lyzY3FaMgHd13QsbjvGfQcs1WS9k1tJDNSU3hGKqouEpXzwxSSeI
uSeOsAhkcW008HPrKvaTXOW1Js7w3hGcPfrrZRQUvCSRMCeqwWS4ckEDwEYOPnVxbDv+r76wb6CA
cOTqCTz8URZtzgkBufHPEIVCGtr9tB9IzegJq+eam55EAkwnUip28//Efo/jHCF40S79ZbtPSp37
V9f+pHeTgrT/Oo0sDgV2LRESKMwKMMjlYYYA/DjPSeXVmYTipIvG0HKAhDWPDRNS2k1hCn/mffFD
wf0D9MN5cpamRiJppRM8MKO/iFSHyi4FC7bLialqTF2gBtLpO8WpJGD6MD/PGJMRnsT3fCBsrtbM
py+RQsdq1txJM9FfnKnaJkn6b/lAL28QEcLvHHdAMn+klSLNuYX+FQGMre0HIvdKUFr9atkeCeBb
VADvNf3ITU9l72ebORnlov2I1MK8Tl2yp8me0B+EyESJnvxMHtXdz8QP4v9z12UoiorRDBioIntL
J0wb+Oh1+covBgUzn2J84Q9+yovE5Ta9zPbOGRSo8hC+plVj0kC9acOi3WcOur2v/BIfWP2LtpBS
St/f1sPZd8Fgg1o7qswC0f6MhE7CH/FXml5npZIuq+fnv/na1JtAyD4j6WL66VuZAI8VxCAxhnDP
u/KbulardRXr7JqBnlnF6DOfUJ52z/9huP2C36vfybzaSp2QWd0OZts9/NnTmiVjqsUuCb8I18KX
2CVSFJMuJjjIlNxJOKiF771R6sX62dOegsIxcoJU0FhuPUd5ANDaEfGkmun8l5aYiMBy3ZLGQ6b7
Wd7VXyCu2AvSH9atX0c3KgW/fFztvvfNo1X0KLuPdGrLLwN2iwb7S181UJD+2RR439eAzauXXfK6
JnfRMUezPlZIuGFCA4bkrKs1giTIgwVli1hOcL5WsLhLzoA8cMacW4DSZ+35pkg5p7jf9fyUfXN5
DK5gth3fq31VAxyvuLFzyXL1FC5cwZZygHtDznGD2S9CDbGx1bxjyxGV5q/0qb1rw266dJBd+9uC
V5dPg2b36ndhncBc4S+sxIFzDvFHJmcQPuT6WrxlZj6TrjHaTRdOyc42kO2TrtpbsWuXeT+Zxfp1
mnJiixTrXhPz5aGMWjbNA0GwJE5N7kJ1vdVXI6J54Dz6US51usHgALQG2NAlh3/LgI+j6DcFg7Dn
ts3FzYZqOfJNtQd0Q2YAXyeVa+zU0Ia+YiWt6Y4jW1I6wqCU9XT2foKDu0bkkw6fn33ILOAKikAu
ATniN+1RoRu/8zQBD1Cl8m0tokTxQk5Y8WDmrHjrd4kAMWK6DGQ04bIZijxOz5vnfXwRujdHvBUJ
7ZQ9W1lC1kDBhtZM1Wp5/UL5+aNJpCChjtO2A1/GyG54jGVS2l2ABX+N0xmWjD9gfQyQ46D3Sdv2
OFsganmiSNwch2Z5Wu8xIn+OVbcPyAd3PnWPpz1b4v0XPwLz8m3Z8kaWPj11xrc4cEtW9Md+f5af
at89GzP0h9mCBQSw372YBFs6Iup0LHQTH5299lpnwZ7adSx6+DSLJcQVmzzE453U0MwKyb9uBqlX
yuvI+kC0BZmswJ+ZMMnsj8HpBd8z8OhYq5EdkowhhCsS7Ypw4kt2tgbcJratqr7mjF+9xk3NGz0s
n+OaqNx2BJkX+EKi/qDgtVvQB6BofWiP4a+Z8z5XF6FmZPesu3AhXnTIGsqTU4d2x4v/HGa7mKJh
Gw5gqjSblvmigFeVhwaIBWP6QWFrrWxEvQhkCPt/f4USqrQWSlkeRBksrmpYHltEzzbWQXG6icIW
ppgC13AQIbkcoSlxNeQ3d99p6vtt1ZDIPKlq3oy0FsJPh6aGbZfw2J/8IOt+QnSjDc+dgZxyMwO1
MlAqtyzP5Pao6iM9dlsUq7T3Exr4quCBmpsiMyPcoJPOZWtLSLduln/N8l4Afq08rdGSu/+n04sP
J500dbnJIfvyF/RwcRBKN30zPxAABdPu76Bfuc7aJVYtdIaC7lidWxY3UY+9zF/uOLYNP6Jjvc3Q
VDH/Ypko5BrglWY1cB34i1//206fIpdESSBYMZHNd81v/gZx1L/5lkHlTcw1kS6EI0NlHbegsrHb
CWME75jmegYOyebVFJDi7wocB9Cl9nc60pcE3OormF9hiSqMaa/ygugqAyAPpgNWCi+wuK5pA1wx
cUTrGWBuAc4lAkkw5U9PYAfT2thB+6HCxdEU2xmaA9I6tzf5LRy3pMnsusFoqZky2GmdAWUvbYwD
zJNFODtK8+zSSdVnNXa12+/E1CFzsaujs0VO35uDYEBy3458T4Qdwc3o5mDyq8Ixgablff/GfS7n
3ul/PRzOxVKYHmn0gD8BJy1rWjy5MbJvQkxSrJvgpvNl6ANR9+hXiFFgJA31srWWyN2C9lwn6SCy
b1MzB4gKXZaeMPtD+2GJ1+DBNncW3u4qO0b0sB0fyPn1RZYCKrWB5cHC1541cUERoGfab9U7RFL+
nEO/PQHGiBBlW2g9lGoNbZ8pRkEzITZ0LZ/3Rh7Elg2Rosu7uhRpEvFzBD4g0dzmK6IadQZEkhsW
zdbZn4j29KACdy3UXPEHczkZR4KTNiY2r6vnJdjkYlhq28Du/kaGjDWXAvKFj67SdCTe/MClQs8b
+ZV1MSc477qNUow3cfe0zbs/5HQwb2UXgdCTlRV5EksJVGo7tbqv9tSnrjptB9IAgwJsKiM1A3Dm
FTk4bw4UA+GAloQLVSJYGZZHpkvXW7QAY39Bih9t+R5BnZDgEDupE9x0vgAmzcUiXZ8Fiyq7MrfR
LACCQoytcRerS7x9eyK96FZraLzX9t95UbfbZVndeGVAiqTOHrJVSc3GoxzBGqueUs9inwbaPM0Y
su7cMoe0Ab9uYvYQ9Oc5lZVb0VqXDb3aS1k6+BU/CE9vPnn68zRvB449WeQPPo6mky8vFRdNZBSX
dvYeJ+N3l4V8J2SrQ8nYp7J6fOwXsjll5kkVQfxRAucZBW0AK/KMhKEs3oKkkvoameFBgjI6OpQ4
1tiGucELu09uoPfTb3P6G8Upe7jow4MjYXuHbQpP9CAKoNPFQPplsjn2nXdIfeDdproUs/P8GJ5t
bxFAy0YzvNQp6GUQK7VW70uEXmZ+Akwfxe918Wiu+4xaUuktyJk8V/DUU0OQaKnFHjBobAgdg2G2
WChiFEZv9mFmaO0JhT0cAeMElQTc8H4aadI742yB8XtHsi07Ol79JYekkmJaYiR2/yTYuMmykBYR
UXWx0DAcQcpTMsyjkbbyykE219Dig/dWFxpbMMGcqWkb/aBBhV+mWp9OXt794PXSwF44tvrCXJXh
nnLj7vxVaZNnbfEsmphayxZRJOTA8I+u+RbrDU9J2PJfP+gnculIVhlvsGBh/KIWwu7MO3oPPJ6L
Xy68q3XAncLBrpipjmhlDVT7v2N0WlQfEqurN/4rYu+v2+AS9H+oMT+DXJL6ZqCdUS+sPt+7OjN4
StdpJGB0S2NqIx2BVbtqvoGwa2uJng7ppaTB/mMJMQo2sUf3tJDNr7ZX+HLdT8lhB+ZrS3ZqMdD4
cpnhIvC6m2EosO0nSHjKrYHS0patLBDLbREdn6bcDNOVmLUQkQhv7zEHgno75MF2epeJkvPCPJ8B
IF1zO1svXPYOsiHqWYN7Egy2v0JrdZtFO4AYv0nHCxxXH0IlRcDdfMGI1YZFtgNrJ9hIoXtJo1zq
hOAjgdsAuQo3uCOo+sTgx6Tv1eBEDnfdUl4XQkkyQliTUcmscOt4j1M+2lwNlX2IEYxojhGJ9rNJ
dOd3BI+0QVjlOdnVvknB/0eOoVMB1Izf8aL58jgMWfVxUEsdv62ef0QGYj1fOx37xgXmYEQiey86
xftJi1sqt+zcurC+5SRPUgLRbEgw5WaMKwYfkWOlY+nHvwgXhCpx0ksctS3jN3iXtP8MfmWy+A1o
K07CLkm0/OqjVZE/SRUacueQ3LI8UkcTiZuWJ+wGYrPB58wgI2HY05VsXxwSH8sbVKgstjp2WU56
SxIPbY/O4Ju6sZ0zcVOd9J0LYVMmIRNfxRpgYsvS03Kymty+kBbxWhPFgsXGELTBuUO8O+pS9ugZ
MXkxWbepUaCw00nj015z7v3+lsZoZGofensdUoYnVP1pvrXGNlZif8OtSkLeTFqyRCl6rOzGRR2T
mZozeXh6TUe/a3ZdQODRp17m9xe4AN9jWRD8vx1qA5AyuNKlcC/RYyR/G27qpoT4awmh4ZY9K04l
QqfDbOZeSaN7NAM+k/jPFe9KlqIHqvBi3WI/TacrZ9aL07k9I2gpe1slHFVAAK1BYbsZasiqlt0s
Fu6AiY/ISym2lVnuckzQLHo3zeO2Ttp+xVzAA2VhqwUOenm6qZkIzT1pSKLVIxDl3QCN5VrWpWGM
N8hzUpgCSHJXgwEPowbYse2Z/aRiqWMleheFAF2C9N+W7O8ESV8p+PCxh7B3co7CC9l1hg6VNWTh
Ppv+hynTYtiG1iH1zMQegyM4hbhH3Xmfa/Iyhix94reqAFzayA/i4pMyBFYr2H4qFlYLHQD8nzZj
WTNEa++SleNYpXDRFpEZJyUXf1SFgg7utYHJt9xqmkUF2KAzhq65D+2cJbHc+V4cvIn5fVWBP7r4
U2nml/7gNXjJgbbhhEOsTq8fU2S09lUoUavsUR5h6WO7LESNrPBktV2BJnTkt+Cl2P5M/gfBVMoH
uiOgc5RBMSJ75G0Ql6Wa3UzBB+er6PxJWWNRGkE86Fby2/pQIZz+Y6+6Cd+7zZAiioGYg20Jhw0m
AmvNLaBV8HpzilHXAC3OYz5NqX8B4BUdyzCpUxzH3JvVe2bLT2Ibxug72PTNCdEexwSxn5TAVcBj
puhiI95XjVCZwfcctFrENQEl72wgYFqA0EH8ZS5DfaVDbXP9m7YvZDMIiGNfp+ryo8tzVCGvdoqo
eZuJ3VQjXvsodphLdJEDs42xF5Unn6Qtoi2SdLzzGnH6ZXY6v7C9aJXo9RWk7RiCFChdplgkPUyF
AlfmI1rwYGCdbr1fxv6Msnpkqub7GGCX0/4Mk/8MM+AerjEkw6sxx4qiMiSls/2RdIOLq3tELXKN
JUKk0hpIVhPSoam4y7LVNdpai5rwoK0Nq5Zj4PcEfy5ldwvRwfaRMgahFBr+GjSqMLdWDpOpaTf/
4To1/EBnzDVUQfiOjp0shDrYxPVlG7HYqf3bmN+6qzOBFNA9Hg+InAqE1XY1tsm6tZ7lZVWLVzJO
InghZif76op6ZnTh1EaKKehQHzPLrh9SK3vG1Es2+XTC/+aEahp1Tw3clU93yU5Z++z2vc5x1hcR
cI0b2wofOOqjY1ZRi3N6F0/7hKYc0y7HcBNb3z3YKi6sJ1esHJYjDN/Z47EGkc7ZS9/CRe8c6Q3g
X4oPNCUtLZyP5xmvz6CO7doIpDe/HtFeLV8KzS2f3lh17oMCKNqIRdqwAg0y+yl4wWShS+066UkR
5nsUZ0w0mxSuXINcudXNigJndotYO8Ow25tks139Tt32b9E71rN7vtLd8uY+zj8UKp5sckumXSSA
iY64qzP2VF5D/3IEPgFjsA9YK+2Z1BJVeh25KfFGwGqhpm6x8qbeJlwlTKe0OHowQb6XVfpN3YFy
YOuCGbTtP6AG/Hn6cwQFQU+HbaFOem/T8OaYUDeOvZmfBvgifcUbEd+3pjVQtphcNg8C3B8gYLKm
doBeN+BV1txKlNseRr4C6pAG+ePXd713ZEo8j6JdhtNaUTU2q59LuY9x4SgVXeQFHOt67IktemJs
6UYIARhGzs1Q3AtuCSs7gavydbRFoDbBXyMusnOjuCnqi8CoQd7uF4emhrUtQgvXgm3j8AH+ijyW
Zx+emF25guSRUduGOGMM5GUD+lstmr0MkGJ7PyMRAp14vAOt3zYfFPc79kDUgkgtiQ/SiODVroo6
ZC5Cp7mTI1Z1nPhZEVSPBickOqnyoGtDo95D/ZF/aRwm62lBTGkJ6QzGYaoUCeOdnUfhcmjQcyzM
i/HpmHfHVZzDynZHdYUcKeSgx0Y5lz89C9mBXaHVbKAIQbaIdfPkwUqOMG8o8VX0FioX92zniWY4
o0wyapVEaa33hEIWPEqgkxXVTgNzppd8FZ8JRCay5vBD2XMKhkwZuMkju+eBLSxKZwLkA1bMl4qf
V13JzKERXEXpzrp2/Zup9BUwJgFl+Ri7tDbXUW/hqJlXvOzO8/X9VtOxovjx7Zn2bnlmm3pUcD2Y
D9U/7nUkAI8Vvb3VWpSYTgZ2XmQ7qd2SLpxRI5aDvgk5+vy1Z1w8LBsag66eMg4CWu2Ric5Rsxum
w5xVnPnGnHcsRpf2FsaGoLf8tgb4vuvXfzx6KRoz8BYaepZi4NkHDQSajvW2vMjF7Qj/fV9eFsjW
ed2t9zfgE7okuxx1lJNKzxf9OtGQEuVKUe3nDTU7mMS2OINFqOGVfIwJ14gwmJyAbYrWTeHjSMsu
o71yFDUehaBHNF0F5hUh5VNxkMdXOOwY4upA/VF47T0DAj5UtXDKUNXg8S246Xt7WYWjGpbvKbOe
15S0Y2hfWQz5jOrJbdEX2stWPNicp93REdIxaBa1oIDkqbR0XdfwYWO92fvP4ksPxEoQ2ULCF8kX
Dmt7QG40Eg/UheyT3poRD29u1w/s8BHRqtdrsxUy+W/katetmmS2ki73Xsvp7P86drRPbsMjZZzD
Dag/ufY7Ar7KZjdEfSjlL5GLiZlrlKVo7R0hFBGmaVg4A1DqvoYUHXpIauEjXY18rruRC3Z75eGF
TpKRaMDrUjQb4Kd405+IBwB7L5fg/JFdKkTBLwJ5nV96iBCnVqMwgNxm/D+DEWWXZ2ok9eiouCuI
4KXo/t/n3nI/Ff/r9Yuob698EVd1YNY1S0WxavthgdAwzkwYXyrYh8J0IP6ba8wjfS2QrsJ7XUpD
VxlUAvM1iorjPhxEUQpeg2WsJuQB3uVMa0hVLo90ttYGbWa2cnNbdbALHu7bJ0mdex0PeGU9yQkH
RJE6GcrhZf3fDbyYC27hZEC9FdTwoGUkPM1MMdQXgQuzZCLwNMH5Ax/cAf1smqKt9bsphW9z+7s4
4nJV2ALCI3hH5M7eRw5uaVA72ZU/6btI8xEh8sx1IMQ97cxDD/hoOUFmu5KL8EWWvM6EsXFCQ0w4
JQ2YwZU6GoiyhW/xjZ+U6aCLZ1p8hhC9F/f8T4eR5UyfaYeNSel0/XgNI1TRgfVxdaDGTxtdyt/A
9HC6R5iib3U5NI1ANITWXOwjrvS1x+3xYoTBYCSU8DLW/SQWlMMFyDDhakK6Iq52lhfJ0eFll+hK
DCkrkXZx9xTD68LZQ/B6QjxRvNJQxT0435Sp1ws4dp2zAmFUMZix4kgYHL7lDPuT0czWhnr0RyPd
KfYcKBUcBWNTKiExYu6l+MV97nrrmjTAAv5tN3PWZgM+kzJBLjyeRZPsliV1iaPTms5yU4x2JxjI
DBsg17zgUZv9BCxsE5MTwWaD137B2w8lKpqBK/WwVNWbc02vKUCCsfXo4M4sAgTbZUVUsxeZjWCF
BMOvNimkElZrkknQweLfO4/rp4J4IZkqnx4v+VkNKJe7clVq6cwTPA5tsbaOfGnev8IqnFznex6q
RzaVTAuRdimpFwqTyo8YPqhPnCK4Hwbwyq1plAx0Ai9Gjx6i2HqMGKgP+zp3U43h7ckyDlXorB2R
usZDG4+4bSfl4nWwlSIEnZ62yPOmt1AJTZ3q0S82rKobyTSAMaIo935MsVmNME//MhctfVRIqJwE
HaZsUGXuJm/+zY2WvMWsZfY+y8Fyispav+oOZ5yus4H/SCBCOIrBHCXNvqQfTb/IwWtt8QOxqIDL
p78clM2+/dat4LU7aXJxx8ymEoxF9SubjuomlTIswkIxnpeiTM2OkNYy1a34ApA9qxMl0slBSxCt
VBWjVUeIbY+nj8wdIHA6xMLOhwvRoBYllHGmrjcIhAmyglq9cHpXHR7IYdPiuVZasb10p3RrTPx4
20YN9556DDnlats8i78KPcV4tTA/Wz4FKWEjA7+cFVfk1XUBfW1EnR5O4QfAJwVFg2GsWc7jx0tV
sbkjWPDmofzwxVVZFK+BwoIqYk2UlMjxuwWc0y6Hv6hyseLjxz6asRxpEPwf54KtXhmilUwyIpZd
7+ncl84Lvn0SgzspA8GiMrX6NAvftpzHQBAhYkNOW9hQin9dyO/gEU2tOHch5fwIcSOZ2gYyjxa5
XSsosf2fCjiJFE5qNXact33G1Yx4VizI7xIrBwlacWJI0ZELw7cwmEAQpGwMqiIgCyuEKpWcdeXn
N/fdTYfXEgFkOHD82+U8kalCUT/BMW7rwe0FtbOQUG6tlemIPBq89rVWK7HMYVGttW87B2cgz2sT
58QqkZYbpZw6e43c8xhaLtUl1OIl9TphDOhfkf1Q1TKHeE9bJ2IB246/epc0lMKQ4fS31Reygu1H
l5EGAM5Ue6Xvefmuf5Asa35eNKno0Cumldm1bk0h2U24HLKLm42OWdxoQ3UaxTIiNjXwdho4iR+6
nnjGUwOfdgUQTcBpdT/fDRfh2Yg3w0t1I9VL4I5mfTA5ZFh68wz/Csj3vkZDijAOCplydc1ujfyz
yQRGiF0zZ+hGbwgr6+fy44OR3G7bVH9FCnpmRnXgtZHdnnEVNZOLRIut0UAiO8KFdZzES3mImr1/
Do6qMTPa4B6PfrTYtgr8FqTixBV0KjBSkeEcFTQMYrEIaLZAoOthIRk4nuDl7zTQzPcs1RinT+uX
dwy0sLhEoH0ohjMuINo6BMIqeDRQ3Zot7YrjEj2D1PEK1z9DF0Odsghre9uYMJjFNtFmx4N3ATbb
TjlwjMK2v4q/wHtOujrpXtGoxx94i54vxg8zqft3L+PLnqHri0WNkd4s5amwiKZBGip6DZJZqq0l
kMLh1qMCZ9zDFs/b8SkTwV4bKt2Qp7w0YFNWDPEIQweoNfGbcAXYvoWCZJKQOjpirgGKIuX6IGoh
VPePCrIGsJ3jaTRiJ1D+3OsiSLGuomIzavnrq1iuSW0SD28NfuAbEuSodwcRv2bH5JBGdf4qnLsy
kToAMbQM2h6pT2K6+rDZlfAH84SejZ/86wz60+3EwzyE80k18Sq8cq0DsTU30wmhvI6EsyA3j19b
oEjmT0nl2yjlT+8XULb8Iw9PogSc2kjJmusWzzt4RdypKcANT7/EqOoH7+ZVzy0Ac0iBb1fW3xho
neuP+I8+otPZ62xam/v8bpoYrrgcaIF+Wk6j/ikOkiuJ/sr775hNJVwpMCIGRi+2NpK0kb8yeDBJ
YLjdOGsNYoM1Aq7q5Pss77djUcFKOKkka25+7HsiHP70IZslX2CEZuFleHyvseJNDXjTOD0DPU5X
QjaiCTePaj4UIhjQXUd9G7NAJAk0ddO2cr2JVsmcp1eT+xLLhQcwOJo0C73BuCAl6xemgli+P0Pf
CJOp8C++WCTtIFBYXvSYgs617WJ5rWN0wYe4nZXY5crnc6f0wIwIF121ODDzxqCrdicXoE8F+c4X
Vs2YyH5yUDg3BuNo1Sic+PsEkNiRndeG4gSu0bJZxr29TZz9hCKkrochYVaUNoS5o/IAPKL1U6WJ
Kj6SKP5ajuEIsgXVK7P+NMKLb33Hbq5kfHT9zdd/GHRCAgo7PTBUTdA/D9JR3Q/hevis0XBq0nsV
Ct+PaAE7BG9rxYKio1yh+otf1sf6AF4WhGJCjolGbuyYcfpMOP9Um2703yh3qbXQ0BNNBHVUY2xz
JBYfdxVf4RR2fLaix1pTs0cTmDAGYnwoNW/Afe3iYwgYZtU2+vLQSMEO9izdXRl+sG1DiY+v86LE
R+BpNOJbr/EK2KHJ01W3xsdDxM9+CQ8PTpAwn86HM3HIjrYswCNk0vjxwaYIbRBMj0B1WGzGvpR1
js3cWVg2rLvoEE/QV6tffqLiqQu9ceK25vzrFcMYYJlT/KIKJCToQXLqIkJ82x8f6y5RPO3XIqG+
yPpiXz02Z+Fsv+GjJshHvkaDOyuRezHq9CMkMAd7aEdVvM45Sne/bSbcj9xwb+7XbG8W/kP88Yoz
eN7Wn50CKpRR1QducNTKClFMrl1iuVo91RBMyKIBxAUXIkF9OvjXYbEYNqCV8wfTscycK3BCcsoE
gwMSjqIZ8Mo5bBZOKl6gh6fbQocc40uQytIuEqXbWwLVMGRjPlmcJ08MSAlXThS3HIBMmaKRpVQT
kjKw3+cNUBUe6ziIqOgPRnvoOzwYLH6uo8VAEtqDn+qDDgE7p2leTByjN8RzgW50XI7waV7LZvm4
F8yAOKa3iLByCNpzynh1VfHKjE5Xfk7foht6S5zitU83dbdn9qUCJ5xZdw2ouUkDBaeHAsVILOQp
UezTnjNPLz9hxja1G77RVmeNLDCKoAYoNC5InQ7Ogct05l7GzLXDaaUMaF2Ix45TtH1f3ZXwAOQe
9fR9k7ZySvkk+gO/yO7wuC7eirjETfUgLonMrH8F/p6ThdxyDwz2jSeKK22mpIuaBNCaUauJPDFA
ky29lt37sUGixM56Bp6SqTvLeFRNq1z8bsB+bZSOwv+/zGbawAxxtdWnyA+8IM60zP0GPNneMcey
z2I3Uv85PWio3te2Abdpb8VtPKHrsrNbaKBaaj2bW2YLRUmW/B8yh5RJHxkoe0LmNOidTjgfjLnk
VzoUUT30cmLNBh3ZVw9GpemUSRGgxxJY1oCytNVPpghIi3CU4Iuhh5aPaqJrS1ZKPYANJKfEG7I1
bvVyxP2szQi3n4iQibNpyaGzFFgkB1ya5lrnGrE2LJ0yhdx8wUIgSQWh3vV53EjddwFUTXFyjldE
Vw/90VcluK3Li/1Z6fCFpFZRSMhbZSju/bYXOztTLMVuspkCsCsrGm0my9QoRGSEjLh7bt8xNsG6
5vtkszn2qVXShi9W/gT6LZuOt7k1HpEjsDQJezd9B1/uTKHk3zFJ1i3c5GX+SC09bRw1kQxBkKt0
wnm1knoZmuGhsNTwDmtpGeS64dwDrhV4flwm1P4X6YCPwJvXqoRI+VOMzWrTtyQpCdlleztcxV/x
Gi4GYa4uw/B2Nj6BhParAOR+QVP/DJR+urUxbbkyBQYtW56QrKczxyoCI0JWtW6LPlfBdqJGe2BG
i9/Lq+MWHMhB0dsm9zWofVKJwlJUg9jPEWAlC9qBWghjKKNX+A+82am5hupooG8FUFtCEL2Zo7/i
5lW6ijOH6jOVi3Uy0D4eIIMUYwVu2JPEFB2GSYHKoUI5I/K/9M59bhk7FfmjpE/KLlUA6ZF2snER
1oxQI5395s5cuj3WLqklymhfwgicveevPylmbYZ0EqvIZ5qjUSfoJgHZmN/ZcYuXjpKDCykLIViY
555wyCgdzd5w4ZxDfEUdwDZDmYY1kpXcrrQH5iAWJEQVNlGhU8+OUvcZvK3g4MnoEfQriY+hh0yb
CIwPpER7FR6NDteLA3c6Y7B/HiBJpYeg6UXZqRdu7Xvk43fADEgR5be7wT2s5mC6hsZKXpMxtLWD
TfU51Q2NQi7pMEs9LohOHjUvYUOGNv0ouzsQUm++860xwoQjVO5hG5/lGJNgvvK6kddyIU/RLw8H
IS0zIfWJqSlnAebk2ghCtqTz36wxGX3HZrQ0cDrV6kRhSDF4TwrQxH/sHmOaHaM7yBPW3hNsYbOi
+QUUksv1jTGTVfo19d+UiP0kTw15V2QYzt8ebEtUiblo3NusYt5OCXxYs0o9oMVDg2BUSnSl4FEp
2VPatVPAIVKISw9QVqCvj0gbI8SdvpPwwpg6EJTabitQxISWqLD3dTu1f4UEbe4QxLwTc54b/l2G
1sdtJxMUePrAT0DUi+aIeNjGUyPYgJwYSto54vD6RJMfSG8YvstB1icoa9LpNeUVskYBCEJVXX1Q
AgwggR575e3hU8sFJz8/201HbTsP+pECSSCtl8Frz7c6a009OgCMGm1AW/juWEYn26oZzcH1qsSz
fT3DUBE5iXcmlt5de6WoL42g0nS957VB9QRnBeIGXy7wya4BNdwEd5dqjpzX6GwJFkaqqYjoraH7
vgeudGE5Tqc4Pm54U1j7ajiwscAANK6113fdxSKqxavFscbytFO/KSUDaWkEDQ4oeKYYLT1+8CRN
aieSZr+0pi2lObH/mryhUv81I+NwIT6F0CoPcngw/IjVXax7+6yDvMuslU9kwOzZEzpR4CsdyAC8
UMeVux4ojWbLY2eaI884wJOrPlj+14ujxwi94YltT5CuX0e5OJBBf1ON5cR85VVBQ7y7Iqm79ne0
v2q9zyx0U4sK+2U12PZv/QRJzSOhMMWWqbDAq9Plp2lWxQgCtvUToXu4K/Lu082DvHrm+BoROeD4
9hA8dGZFaeGBKAa1/JZIvDAh1XAge4duHYdDp3zAvyi76wHasyGzaMEsp02OdAgKyItiAUQN5jda
K2ltymNZ5Dhb3eWro3Vv1rh6ReNmODODAzQGkfBpNEckxDwOdA+hZR9/lHTjaj6t1nw2rXn/XiAb
c+4HLgLqaAfGgOazvD4L3ZMOFkXa9g5FvvZuuG8tL9erPSwLxeoYV38symCjzcouuh3OZR46omx0
5Ohm6foJtqQCF4MBh52hPMVADYwS6Z87/uX5JtsNRZX6qapEOVczGKL/2wOzjPCp2KQ7LQ2N/kRD
aIh04pymkOYdmp6xPgijLgF4bVNyzuCYSqgVhscrlOAYJEdIF25qwQzSM2RquQCBGds/VRGyGXHE
XPStUWX1R3A6BXIAk7oprhapyhaNYnpo1mIpK9ZmdLmBsr+BvGpmTdTRnE4u0o59fTdojT2vwtbr
NpqRZIwxZ09wzEZxfAw3VLLnG3jFa9IAaB17xQAbvPrhN3rtbpqIwZohK32p39EEkweGJLXpetob
rQLQsCFtOb6w0puoPh7eDxZXvfkHUisnDnsrm+mgCyBOHUpOwLnSJGi3jVtnO/M3358AYhGrfDFF
2NEzczUTVIL7UxxJ0+Iq7iOAfS1J5GF67pxR6XCHA20NDKmdMzwtfGlzslwrgSCpmQ52rcvFbitM
sRCeegfWKc3etDfhJNm4o/Iaxaok20UTOxiwYw8i1CpmyVCPosIr243erNqNMr61O3SuQWyUU8E5
aHykYEcrSVcyRrwTBS2xfsGIjRnX46IRukvqQcOajrBqd56lGq+DNOfBBhIOKEOPs4y28ROM3Udn
oW5+S4CCu2EnJdud/i4PBgaYEwmBouAM3hPpg6fLv5E3D4qDgm8irwUfSRX5U9/MjvAYMDAVFNuX
8ojWoqWIIgtcgOpjkpisFHoq2S3/M+4kQqO0Y9dJdB+rzf0aILjskZfvsPirFd/OyH9yfSvC+96W
Sc/j0F3CsvC9QOULsXH4/lAo+iwduEabCyoWlOGdqB5rMEgc2Z7uJhpjKuX/OrTslbtYR+A3PHwa
9/hIxbYNeNXYSRsX7EFG96qlgGpq8S4urkS5ZlVMo6xIaLtr7jO1YBlZ7DOsgSRc1pkds40Q9FBR
ihQcgtMggsuv8mtfCFhk2CkSFFn6AYYTGJPlwOIhdl49aMF9C6L5Qevyh3zpedQ68pDGrDKdwgrI
CwbPWBRyKuuwc+DhH3mqtaChWGDxopowym+DI45yrkhG3AMKTyx75WEew3+TkqMXF1JV059O357T
4UrL1JeXiDxH9GTNRkrQ049ymrA1JwU6YrJlupxYbCkhpkAutfK7Dr8U2IdfxT6gUv4gpHEvGr8j
We5IusOSL64KsUEuoUdcJ4MzUGvsirLZg51I8rzq8hwJoAYAALcwNzvcYbstHOpwxrTgEAsQAI1D
jJIjGxvlMQteZDv9Qa0++kAgALRNnvbSFIJslmV5Ns4MhdXJbC/5FAvJIB0D23rO35wF+22Yyy1F
rQ5Cy3jSaGMGWWEXFGTr38hg1ScVk27Xe0YxFIDrxsV1t/+SWlxUnUPpr8/wjkTHmRff1+L8iHly
L540sSZCA7wbWfcDeMqcGuJ/P9V5B/w4u6eJkh8sh+iVJ57GmdbB1xP3XROZziflAgt8PriUGbzO
gKLTV2DD/WKayJUGjX3z0Qo/jDPlAL4yW68+1ngr/99nU85XSYXR2GDG8FxjbMUKBLBf/U0HgOv7
6GvQG9piUzNrdZx2Wmuvt1EatZO3vv98SK2NMTMdG/Eq3FERuqDoTIZ+TLfgMn7p7KxmQDAW4ir0
0uOwG22FpHc2YQ61rBtUFmspB1OiUs8+YN2JIyy3x+AGCn1Eb7gIA4Bf0zmz5nU8dZjl3NtMvmPY
vCaZP7QpG+t97vscicwjXj+EtvhNexsWSUvOTepAxd32P3kX+WN9vA670uUA76s7bFXOMjuIl4Yx
wpToF6TLVUhl7sJOmUP6I4zbYhuh99D85u3uro4aj9zCHq/ulBC7TKk1d5/A5KlMgTFt1Qn/VYJF
TNKY7MsbznD2MqAZc4d0sw362bp1r8QwKL4NFlvWys7dAo3e7DLrAMf/6fsdouAOlXBJj0kopog2
5mMm2uNQJsRsgiFbCHT37kKr3lZT0IVlrvrZfV1kolwaKbQArrm8gsCLjmsoWO2MMrTmoE525X4+
oUJdxQPgVKjYZmhnC2wHeKzxTlq5DL3TDOH8Ok8xLqXBtEu1DMs4l3mGqPK4lpGuFp3HSm5BNb/l
PDfrCIJrOl6XEeTA+IcfIluxdQGjJ+oVvY0BYQ85D+JegScvjG1QOKti1/guX7uzBdq8AOmol6uO
jXVJ/J8oZ+ImcG1BjCIJO7cjLO/loSLRdv1WdeCa37IxyphMy/EaOI354/L4TAdCzgZeWVQdKQ1M
31ztkuKIShJ+8hfXjTMdmsbpdH2kVE5VtjHJ3QnKvwEayA0V8MHwiqKCOzusXbKUT3NYQP12eXiv
zvGnelXeyoDpW1ONMXvjp3AtQYeQGax1XKQsQAy/21wGzMWVNsSNbAc/bfL9uQLwjQdSaw5YZuW1
i5jRVcq5oi6o0/WGm2wfeI6ymUkHjrF7IEDtzMZSYD3Y9jmatAYa0tbbKxwRWXXbEc1Jcoy9t0he
BHxkcZwO3xeA8csOjFgrCUBJonOUzV16BRx06JqnTfbNELvSAKu/OSL/PlFs8iBUpL7bOnQzc8Zi
DTVzqD8h+sEAxaeDAus0rTfpdn4dJEwtfV04OqavXBG/PMtcVI2MDzUgRgQrqEuZRTsRWW1sEAce
PoCIQiPVLqKA2NRRNbizSVLWcrUe5PrEyeqqro/j4ESHN+30tRPsORNszO+XOZr7/Nj67CI4nmCw
IDcR7oIOnS6dlCKxFckRWbvmqr5DIjAlCO2AN9R2mEmcvFXAjSIGzG5llsC7BsuXa3lJv5v8tlKx
SvdFmeyYERK04kaiTHOMSv3eaNYym4OQ09R9dc4h2uKQKu85e8vZoLTNpYgSHLEgNefVgoIwq+nF
NnniM1ilaQR3mWOcOnVCSc43851s5Xew0AlwmNEPUoC1cBd3Cw2LP7GAGefJWOVw9yqQ+66wKfxo
UDy3OJCiSwx2DGjR98IlPoPA83+vvSiUrYJJtQzzUIlAqutcu65lPYOSA8QKQUS6tofvUWHg0Fuy
ABvcGqW/LYmQj8JGUYk9YvzFY+FTPSdNdNM/e8BGt2uGz//4zVPpu+NPoqhxuh6iAmnPWQr3eHx3
oxySDKLo1z4UXQDHcNbHgwQD3k/boHzt7B3qJE8eRzl/x76pvuUBghm8T3P9AlKreRAmzre1QHLZ
eUvJs8lozYXqIDmqT0NqRBu+P+q6/Jn9b98k1SyRw39cmRbFz6oiRQftAfSKw/xtLsv6DKBc90Kb
D0/nmpo/ZCfR1rNgzj5BCTbhoePzTMSGL8e2XBl02mW0gjeJiVSE6k8ZsD3zSTl8/oupQO4fh4zS
QI08h1QktNh2VgM+kxpHzHymyTJMx6zddFGdWYWB9Dgq+ng4muqigjjA5j94B28HMBJ48mOXCVCQ
CRPoaJlQD+U1ZBhhwdqIa5T+jqh68u3v9zwTVp9AIWAS+CxxMaboS70Vvda2qMBvNaYDz6kmk4Pc
1KIcwBPKBKpat3JIbwdoB2FJ3tZtIWtPE4adC3s9sye72YHX8aB6h34TUQKkFEDegG6sjsH6O9D0
V9yeuFD/NcWAp46pWC1m9YJ9/AuyayULew+0ch51Xk7Qp8Cm/ZVDz/1zLLbsc5ZlAnQF8bW8/EdQ
GMSlPOIsQo7AwaG+mx5MaGB1ABvFx9KqSyd4DcvsRIJkiDkqfG1S7i+Rr5A+O9NDNHoHkXFW+nFE
6bktJQQBz7kaRBl3mnFByYsvOtGFtq6pxuM/QC6rJNe/OmSkotK+c85DtX4PtEAK1hffCSDMKI7k
RTTFtY+3s5Grc+TPbNs8XNA52MzVh4uEWqY4Z7fR9E1JvaqD6MsMbcFKeRS0Di/cqYm1Zd/t6DEk
6fkqiaVPMY4MVEW+IeSs/yVjn1P7NWPYu+MQFn5HUnjxx8AdG0yayAYXIyQ8N/5Yy/rPZ37EiO7Z
uvdT2SeNAPh/Gmp9ZFufKrCGE8JK6dxUk8/5aLjyMHebNaEm9vrg6ZEez4gW6uk837GRzXyzTDFq
vnkfeptro6g5ZaWrnVrLBacs6p30Wt4JECf/f3F5uNy0tmSDJp1tY24QaXD+mAR8gHlvtF5miy/t
FB2I1C7tvhmU2cXy/cLWDjMPwLcgyRPttJGVBXn159BPwxleqoOuF4w7UtVDVgmvcGb1/d4Yi6xB
DbgkdVnm5Whphg6sEO9I+LiU/kS79FimJSwFdAmI9q7T6qRZx+KpuNnmkJ7ucTeQ+6SvrvOet1s/
IRv8IsfVMfgN6/BQvDKIYGU/dTJXimNgu3AlzkgbmAvouVK6g0B2/MXhLyyrnnAObx/laQhffQGK
WJlzIMLVo8e69eIfFTgAwyERS9KEEitX9yfe5n22wn9l3Cx2sizfP+1ty12V4J+9NYgwdNlp1pSB
C29T5aER/Ln344M8kCadgCtGWsNmmD1AuHqRMfA0Vclaa/zrppkSTS6sxudQw+oal94JifPX79+U
YLLcoP1M1vsAAY2khzuOv7VFAM0m0/xeek2JjtaDFKfC16e7es2FXUhN64m5PEnXlIxK3tfsnJDN
TbHYz6RU+JR1TU+OXmdzG4Leh20IyfzZN29vfhQzBFrIuBU8vwspi9yn2wpeHLFKWG31G7l3Va7j
JcU7Me1yRDTO6LF5msEoyTAqia2Y2MyJW7Zkhd1duRLaIcHugMTGmHgzMrLF10MiG6NvofxFDii0
EtPYg5v+uP1UeSk5KOR4IDdWSeOyctoXyTw4IoijdNxlGI0XWiKS28Gk5v5XVSBqyzyavvKmIKjW
6JTfVXevDFCEiloiT3aEJ06TxjkWF5tNbN1smg37zmgBloDCQxPQeOLyAcVTgqzjTcfofo3SO7Cu
xDMGBlyIOMJrsYWPp/Oe/hB6zbSK554VsDXw7vvMP2qZHNKz9i6M+8bvFAx7686tgOlkoFxS3X3A
Fw8qk/0lb60mIQt3kdE+D8gs553RcanP0sU9ywGuYejeUkUrCngTfDLLDFTuvle9ZpIokNQOfd4F
yMn8WnZZWcQ0KNXaBthjZ8/EuHVXvS28ZzUJ2tZQYT+uCpoF2aWbQ41m/wmeoiFb/s5ltZbdXo1e
oFy2S/5A6Ot4GS4LPQBTVIJTbPy5MZyhUPY2eYDn8v58h5bKjdoqj0dZpmIWurcy3DvOskaqwTrM
1EPk1B3fkonuuL206uWpjIzMbe1pfQnX/vvy9cUuYHLpTVdTLyCPFXC0c+iF2MlWkFzVpvty40bP
U8HKHtvlu436e3OofcM45LC8Q9rI+FCIR1zPqPLJrN34W3OwNW2Hdj/iA1v++TSn1vTy+gs9GJL2
LMZw9XGbIBu5bwhiuG0KgFAAEH/OCHj+SeqryYaWhDI9jwqfbJ/4Odslwp9tnc2RdVVu02DF6rXL
ihu9Fu/QxEiyUwbIJ1d3Oz2TzHlMddgKCp2asU72pwQzb672ihwmDT3voXfhJdNzy3SRICSF+nV1
x0A/kWcJaTp8gnxRduLXzLDlSTvBbaKRtbY9dHhOBKMmDwIAvPGX8FoWyTR8chCcZy/Jh5KNUiYg
65FqjWZKD6GWlDiH3yB4Cr5AACGkMNO0zGbDoVgBbl1hS8Nbuk1Drqj9zHUNsT/uPCP1r5zts1Db
ZBtdGVII8nsgx7+T++hp3ysRPQenZi/fyIKwY/nncQ3dtf4fG5ftHdrAImmExB4Kq+XkEeU5Vg72
fSSTFr1sqnRUAd/Wc80MPBY9WWu8+ixWklPb/4eoWCvJFY/OJL40fEGuE1kZR9xl5Q/xym8e2plW
QldHVoXMr2dSxq7gFxVOsppjBty7/iVz7vKvrEc1ZZJqFzGNF5/JMALvfrsXseSswRZbv3RxO7wF
xYqN0a+XeSjVyQPBpFOYqH+mKVrSoygIxnIFGmg9wQHVMJzp0kLWmme3plkyy//bNbU0z319U6kP
vz4l4P59NE7E5ENMZbUc4ZSy+95aV93zOPLsITN+hsm1vaExLtUAuCPuEeHvtMUZi0r1x72YyegP
IPQnrq6dJ41pp0dNlgcXeArgxEtvQs+WF6SwwYmRytZqv7AYxoaV9LmlP3H1qc4f2Q5ijH6/PDuW
npDVINjZ8z8/2i1mhrKs7cVqdDV7/0om5wSBBHagmVoj72YKfmdWrv9XcOrJtWk99tYgV8VmuyCD
t0IgUk6sqoxNd/2Srt18nreHf56WFLPSn+1CndC6DD13E0xdNjgDWcVppMUZxxDG8/YzPFbQDXXU
mE8p9+rNr1QWn15+ay15hEPjYWWzd8bbRTWIrTsQ+SU1r7V+/f9Po+86AzmCoerDkelRa0M6OLgK
xP5U8jEhrQcxgAofdsmPeHAA3Mir6CaqkQTLN4iNLeVXIju1W/H2VGBwtdOiyhPxkp+d+gZ6hlEH
qQ9qRVzVTXo3paCfqkqUV3z/2aVMyhNHRl1fZkRNXkCbGnjD3Ot5scvRbgOjkSHeNtktO7zk65DG
niUWxakxEDD6wtqP2iRqy/kEvbjZNIPhGFpNmt0kox9VlzIcKXU91A4QyiOtcu9kutd+APNjrjRk
eUoz0IsOuGxnv/OfSOE1J70eJ6aFarL3sLb2vgGPUyEXzMoXHivJMdn8B4s8t7Tbs6+EsanjwXHn
qT0zLoazPna4E0zwM10hkg3pdzIRTGDYgvQO9udjr7nc0FINyjIn2gGAeVrlqHBCrpgo0phAekWE
tlB0+iFGY5cVDeNr+NB19ZDEWE9m8U46RfzKFMu4Jr9jGBh0xWHPzu53SuNIfs82FfBxmEsIkUf/
PVbohZUZ2L7VtCRx625JNUz/L753e1tOSVLFBLqDAJWIIu58WgxUsma2Kce+hHptMNpNI9EiBn0x
IJ4AlGIQhz7vZMIKLSDw9EhRE5gGPsZ3P1rmvOgvVGWGgg87+Cxu+3pFWdp8AgHo1jqxxmdkcSme
2kn7xHu7tOoZ/l5x79BxfHFyw5hVftL0hcZEGTuWjb/3nAPommpP4H4pPycpxlrcSGP+7E2cMJtO
AJ9xpMEsWgiwl4gHhL4sKTkFO9SfXfULJVNtMz8IzSlOPMLRinDVILYTT+VnljvpHJj9HsRLmyCu
mVYrju+tEeX92S2kBg8d3Fv0tG7y5CNT/G5GAhnioJw6kr9aWkqvtiRd5hSk556GPzi+gt9PD7Gz
m/ssnibsZhaw0v/RPUOyTM1yOt9xCoXuKybo2bpfPcpfyg9qNhLdeVnCljDg9RlfYxQsK/DzDw59
Pq9SSNjgscRxLCFR6HAXvBLt2L12qmJnp38GKIXYCqWVwYwYP0ZmdHvOYrrdZFDnAW4O/w/cVyNx
IHNL86BHp3XlnObuX9NsI2pM1rC7//kS4Ox2RTLSMgkQ+Jq5/CtlbrPmulUiTdBPx9/9h4rpIDLq
AwvP55VgNOWIZqvSZLk8X2FZuO1+IKP0J3f0Gdp0FsQb3z2Z471/McDtJ4ZVxv6XOrBbRWu6GhJ7
/ZDtnXT+0DS6OBodoeuXsKnJ5SET5TYNJuGqNYsyrQyWQimodCmcpPc0CY0CgXvSWwTPZRkNCezU
PWy5XWOMFoS7j8XTKnuivX6leL9xhKYNxYnNKJAOiMegfxbcRgT0fWchX2XMaCN+ZmhGDeOrLsvI
gfGPsnHvRx8YSxmU6w2ihfi8a3b7hQWa40SEc8XUEJ1oh/4JrByIZ0Kjm9qK7f4qTBZhpLuQc9gD
ag1vOO3IfHPdMsYQAeLCgf1kVzq4lpDOdk0PQwZIs0wLfF/h4vGXW/F6jK4vE1CmpdDkNB8zRNr5
Tki335Kqw+wV2KAdvRgrIOAhe/DHRiwt2WmNjqyINrXzQWUgToywh1ZUHI4VjK0GpjXaMs/8sQK6
17TdQViKnrRMiDf9oy7C7w8zcirlAHm3ti8andjJC8n3mybolMRL0lNnlQuQx0DkP1XYZqt8h3E9
vortUkDUX8x7L/KyCaBFu6XMUHtdoggXSa+39PdZLUxj4tZyRMXTvBlvHToYcjJZP0f5ZOp/r5YG
tvl3GOpO3fcEk4XFnPDrkzAMeQqYVjsH+Rzo/5+WG0s/hzP+x2kTJY3Kpjx7sU1WlsGr7xOoyRpI
SFsRCANHxJOk3+76HJpq2mgG1oqNuDVi/zW1OflurtMD1DSYD1YyoBjBT70J5a6ONx1fq4zqfYmu
xdGzkHfz+PGvf7/6XTEF37O9Slwu6wioN04yIS2dGg6dCa5afdr5hFhDnpfjNM4OhJqViAcpQe7O
UBLG3MtfBrUYPk75+l1cqQY+vrcoSygV5hBD8nNx8woJRDYkZonD+jOeIyg2ZrqDdkZmeUeBIeM9
siotKWxzQJObtPofaF98SDwgAlZx3BHgtyaeqNe1xhKyt3ICKNsPnseOqCjHcN8Wg6PVSv6hSJKJ
OqVqt+rk7f3VoXkNA4Og/I657Fy+ZV60kqaxcgULfz4vY67mdZf8tf1HH3lVOz01PRI7NQafQR3u
LxAXT+K2qz7YIj3xRhRvfHOIGDK+jEggStRTAzVQSf4SPsV89MbHFyZP3paZNcmndnxYx5tWkD98
Wims9zZJH62O9xBuJhuwbJ+zpV6m/Dtelf8AV2551u3Y2CCvu89pwCxjoLPMNGjU/aOAYw9b1Pvo
PBt84OrV6UV9YmGlyQ1zn7soDY0cMvcPAqCMwQWdo8s51sufPhaH/XfIASNXobSq1XBC4bIpPenu
vntdtUx1WxNFPt0pB7DxyQUoS0nDkxVIiy3e8RqMui0Qq+Z3TiNQAJIVBo9Gk0ELYT/ixHgPIxvE
hP1i0ApXUwEfmRkWX6gDUvk17DI0CilXJOuTTB+o7ZXwe62BFGqOiYcrDGBifqZpnqTy/1ipyWHA
2iNkJ69yTd5x6wuq2JHjj9Q8oJCk9q5us/cBoJhzhVdoxjb2n6+RNf8FbZiQJOvxrIVhqvPRvNWa
VcczppbViDX4AgBOuexGY07D42lRYs+MS9ivXKsF+EQTrTnOUXzzKgpz5bLjl564ipwKR8fEZ4Or
bt3oJdhxrMB5+OU/2+xeFXlti1upNrr9AuXZ3eHlTu65HR+SmPVjyGwIYO8muMKatkrkOHFotBwK
7IIS6IO4nzUn183u9H0rEoTyL4omfNU9sskUX6Z/tCbEYvMyLqsYf+jY4cbK/0d1/R7fV0FDuQoh
+ZYaD/8oc00Uporp/DBNZkzhTNZgsdzfUPTPnwvGk2f+UwG8bdjVH40n09J4V9Yd8gIIGrEKvpLd
zQBKOvVIxbDwlc6uliDbU5flrKPWjHDRsbnYsIbl/BSlbn6v6di+e1+5sCO2GIg+JsKNYtXWtazn
/Vi8qe8fLODWnpXlJyCXATz6p3ZjOvp4zf965znerpgaUl/vxZLYhBsxfybvj4xzHdusFl/FnpjG
WRZFWcEWzX6Qw6NfNMOoBWZo5dbya1ptYZruDK5afdBTD/Itori6cAR5rykcbIzHE1BTopTPyKM9
gWLZCqJEVJMBzQRKKERDGG7ZzglC7sDW4ls+y/+S6X7OG8BukuSd6gxX1bjjc9CRDrCD5H2OtzL5
uOHe0u/7OgvUF+YJl6aHRoB2Jo1pZBuISuV1MXsUAHtWhrerH2i/8CV0zozPbpT5SQmsd5K22UQa
hJF3ASiSX9+fZYzaowr2Q7Kg0oKLjmD7D/5ptq4SnSeE3eWXXwMfVU44IsUErFMpJAmDjcth45oy
gmIG+yjnadFpjQs/JXX5hknDSXC7qEdxsvZeWOY0ho4+V3OnfklK9OaS6Y69hVWpTx8Fl7Qf0c1R
tRtvgXV7qw3GCIH1v1cbnvOJE3KKIsEbRctHjR959S8FOQNVVpJKY/g3G52yYvgHNQUtIKoeYfIz
GzRWdbaFmwok5nX3bGcR28O61H46wgg26mBicgJoUeFZIUmwF/vu7XAn//z7AypkfIxaJIPssW05
D+1nnSjPPsukC39xv5bkoESy6LBmf/GUuMynjaOfGd4f02sMNvKn+1mDuQX/DvTcIP3ErXeEwtkh
L0l22fI2fvG92DZyO9dJBn3+Y8OfANpYjOYW2n5gEYlPkNA0nQ9KxcHeShB5XDkAcW7F5TbU5L5P
2ZtRmIdx9gFdsyCmGZWQSmNFqoN4oAlS5XgvfycCT9pYOaHmbFGFEYhVAsafOOLxveGUHY4l/COk
w5ipWpo8a3hvMhF/bJIWA/t2HjiCc0geK43AXXVITgi9+KeJF6G4fTYnQm2vWsVZf/ARsywqSljF
bLqZM6KUSBUDfMv0KOGbXKhAeylHkibfjcN5zaOVFPQVPDQ105OuCJd+x0XlHK9Sq4wFUp00Toe1
nXs5KH/jmhgEwQARMy4dFu3crOmFry1p2pjfFp5z48j7SiULXXMnUkC+te1gcgWdkQ/+aGkEyoKr
RQ8qmI8RqAiwiUUNy5KtrEcMJM/2I1Ymw2jZS0NdCIMHBXh+qrWgF7PCck8PD/yqd/8UuFLZ2h3G
5fB4GA6pqZcK1ayAmxZOgjtKyXZt65RaF568RQvToz39mUY1AP8D968Yivx4O5L/KzL59IMAkS1I
vd5jcgG2XmieeSmkHimO/58Qb+J7XA+JrFBaYKuTE0hfKHRmS/ruMmD49Cyi779KsEivph7j+rJz
RWZ1OpvGzxqNo5R82o5hqLEbOrDinie9D3p/FwiS4W5beyLBdYFwjGLUKJLH3szzrfjVdR2mcyie
F/vLHh6fboPR2++WJCen3/kZW8XPOrUXMtw0CZ+IM2SeiEsbSN6eeX/36Sr2xKKG51UNgfDea7Mn
YO3GHKKqw2ygfZoDCG2iLNd9NHHm8mI+euEd6puZMau64WDnpNEkR7ecfynBbvK0hUsGe5vzX/QF
xNSk/RVEl63Yx900NBY5OrPFWWZUr8gPSI2oKsN+0hNf0kN08+3O/RmQBjA2xHlAYFavZG/ao/t3
yvY/dJ6kbAcBpfJd0pAgaQds6gWQKw2nzokzALELnH0wbrl5laLwugZY9wZKUKwFIOxwMi98S5/7
MuGTt1ZIm1DGV/OWBFSwY2EgCarHBTQbIko8rssPkGdofs4FIFG5u5Yf54eNf3WO/J2n1IxlDheP
NXbyPiOPXlopksKwRTa5F+6NJ4Glu+2yY9isochAyg1vGyuHZhR21hCjcYmbkwJx1ZT8+fIv1v0N
ZRh4s11vWe9GNE9fvPiVLy9vRBuTWg1cYNlk2Im40/JAgcKCk5QfPLWYHwwTSt0rF1Mpnxo0qsJB
Dv0CTL8dfsV/NE912NG9fky5KeAkyuknOAJGGrrRbrKLTTUXwr5gweKf8Q5hpIcAJ74J7Y17rz4v
tzRGlD+1c8ZNokJ23qmG1EXxKszts52dWYw87eDWMzF3H7EKleXRUIfFqttMsfw40KllLof7RBaU
kbza8jN/PkCHpdSrcj2TC5ZwEa/E62LoBR+g5J/8x4+riXZ7DDHLQy04p4sJhl+6vbjrskYnrduU
NKgG7sbDRbZrxL94C85NXlSZKPsL+hSmMsYmMDWHjp4QnrQi8t2TYjvs4UEk03z9mS5XRZ5aZVYz
1ZFWiZy8qO2TmRdmsQU0N6hapVHJavxOK3iyeeTbgQEqn1g22eEc2FT6eJtu86EyucELZrGDkcwN
m9VDhWHka7KK1+md+souvzdwMJ2yPMQcIYZsXz55sBzMoDpyQoAgwWZ8SZZqdmKbbb4bJ5283GZ4
gRcLDBqiwXpG6xIMpYxHDqPnzke0UkxZY5W2HG1wvf3K3Tf9YtVc72CgBvY8HkU8QwHUc9vU9LVg
DzUMXUYbmIvCxtTIy7LVjuhFk7Ow36+Wf5/i0QBR2rDFBZVuEhM7cNOfJTv4NioU3UOOmNM/S4Ce
+VEIWgVihDqFW6esz55pHcMRxtVNoCVLSoeB1O9Z+ZDZliNnWi5N1PXq6+3B6HQx/0RaBDOFbKeS
pHeZXfVKAGIpvcZs3VD//eIDvaZQm7OKd2G56HdpP6ERjaxeZL3ltWTfVLpevJ1h/rLQlQKdxamE
y8il5XN1+3bBVMQfB5m4nCPT4y9u4gLIKxoqoAKMI57WRn1dg/4thF7TPkXJXfXt3Nml59EOBAOx
xX7OjJS6NwdYBNACjQT6kHzU8TefoFXlLHcv1cWKelH18f1TsKHsZ36KMN9a6wz22laUAPX7pkk6
o87A8v44rjzNX28lW/O6D9Fi/a84jhYYJILA8ug8x8jQ3pEtyH8IvrPHGUPs1oZaYko+vxvpR56P
xEs28yWktlqTRFZFHir8GG2LM7wN0jipWqSNDyD6nm03ZF8a+AzMKZQ51guK99x8tqTJacMTDV9k
S00uO0HSJnYYl0p4wxuHs/f+aR7U4QGYTf9xX/PGYwzsYIkdk1HEoNWbYeywtuodL4ebI4S9PWhM
29HHFNbW83XiITdwajg6qAOSZyx+NUz30ShqJtoQCMo5DPTmOgwTMGgBcRje3P0bZ4vdPuU5OXex
ZNn2A/BcD3tuyiG8qPnvVUbyYTjzT0F71aen2t3yvQVfVQnSxIJeDHU3PVP/v9gT7jUGk9a40ytR
OZRWlLsP/+vTWkvBj9+uhRLaVoQRE38Dg9Skuo0eunjl++KViFiuPIcEg0jV4hfDRori2NUrarym
CYwLESKFEHY2bBdwSKSNLSdC/VbF1TB4990bu7kqwMkqfHXEZ3pX5da8uMUu0gpaQRdytufN/Uyl
I4qH+7Eji5mSJ7dWwv0maEgDkXh7vUl5SCwu8tuvn6OnnKDGwRnUUe0f/ZPgyyj0JyI8QDAYbLCj
SfcVZVKcqMBDTupfdprjnlat1lprnQXWli9MfV5yHEzFecE9+eew3cWF6wRN/gJYIvfLdw7IRrob
+YqyUgRa1bcRkvOoLpUzx6ANqlhaxVtF6u3Mf/sZ9OUvq7tyq+3u8XqkrpWc3I3SG3Ea7+rg2swx
j59F7T1OocSBJ9TV+MRaA/vFySjBr1IkHxhrDJGAFieIv/nqaiK4sUThVdA7tD6d1U/wg/xyK8g7
oBIXLKd0iChEesGFqM+7/qkDqizCSDi37O7CynkQjFk6Zp4b1IY4P4MhDbMTE5JRP3gRwxfJ+8fk
oDBRlfd3UzzrGKIuPSgt9eM+2l8FrircJuo0EBA4gVK83vG1cZrIJXXXqRTsTZHK4gs03Yxu30Hk
6VecqhzRRDKf5oTUPic9Acofb73zJR+dCs0hUFhsAFffGRnP8bpDeRh/qzTshUDztI+AHlpJRKOl
wptqmTl07FnAysYKHDm821Mi1j+ZRJpoilqyJ0wvn2EdTEA1Bte/XFn1NDaL4mMp70/nr+PqX4sn
yp2qEUW/KsLqyz6OoKokedK06StnSdkVAFJ4z/WKK/JYmYncGswwPimDgdNsfJpF+vB+lIGk/Azk
9GCJkLnf8eGKWNAixvtCwpPoMbjImx7tzViQXaMqREO8nFsXp1HER7Lasftu4movyRHEdsPbGWWf
POcm9aGezJIhXeWL22fhMUxpDVEAWsUTDW5H+g7OPEJcRRzybG3RGjWyzWr7WqpDfIIxUp7QXF0r
0Jv5SyxT80Y1/wIzTfEp2VAW9LDHo1hy1/is9KTsEjc8QeoB1u9MQa+SDu906k6xjdduH934S4eJ
wrktxFlau7VaayGTXui7MRJrlJVg1UNm/7lI9ExhhZgLssZP8kHY7zUrDMRGHg/eH2W3m5op2n2K
5dquADjwMomDqgPFJjuNxqMJtsEHfr0AO1lssivk6rl/XPWSCLUWcIUM+J69PvcGNgorowYTZ/qx
+FaG5ieFbbc1PDVxugrY2gAITcW4flXtTSsHrH2zvkKdgw4WqMvPlD82GUvHj/5xJotuuYGkOc+n
i6GO/IzFPxWUnw4TuuBlPMQIPHMdzUbdIB57G6+6amdi8PcUfdMRE4un3dqqRPkxwE6n7m5aH8Wv
JeK4QqWLR6rsQ3CoRvL+MkX6GdGCTNENvPVxQm/U52JHAqGbNIfET5rfIPvyT97xoR5qD30JWG72
JeOW37Us0jiOD0Wf/KVJzexPt+7j3cxzdki1nH2nafhU2fpuuHI2+2fLIKIaEkaeseVUEf0qcvJS
qHNLIvvt7JFnGbFGGszqMXXppMQHbit8LpfQ9mQNBeY48OuOQOHiZsSo9s7V8iWmFUfgbFQv5yU2
F0W5syLMLuzpbgs4GqgPgocRQGj6lNRGIWw76sj2i3RJCtjCnwK0rgUjGZSm1ngSFOpMVhQnV+Cy
0cSj/uQ9Ea6wjj3xd/4F4o8jZaj1SLAuiSMg+0bhybNEbZdkqiQCGWXs+lFprpHlk1MibGuyDfxS
rTqt2kEc5wrF6olZGqs0hVYjuRhXKS5Mo57SuHlzC8mZj6l4ofPFbdphVG8J3QVyUrQbZx6vKEal
eQUv+wT6FjQ+qsC/zBO9Tyney6dpgRkZaua3qQuW6LVFWxJE11wHkUjy8YLP47yDiXMuQpiWMojc
lhi2NoAoDn+R7UzkgukayPGphObl6ASgTLbbAD0PHRrzqJ1/cFcEs10E1+TZjoyiIlCiW/zIELaM
OA8ajPnaREPeuLg9Gni/ATSNeSl6VmC5Dd5vw5G2nJ2ohRr7JgCao713uSG+KCZDo5IFC7Ckn59S
8ZBL2GvvCu7eO217Gq/SXWGLAjUl4KvndzoudnVtTUdUDc7L6Fz17fLrksaVj4Ti1Z/THSb+nmGU
1OyLChCQdc95tjB77OpWLorXV2G4l9jcOnJzrLcW40Yc/qj0QuaZ2IBiqXfWmxt55ueDNX/J1GDf
/m68BncohZ+3ss41UM6+BzK7B8eayvRA51z20Fe0a6uPtDxRtixj9PdMyEFe0JE8f92cuEVsyFmW
eZ7G63GiOhRYwXxX5ckqD5kW/FDVFofg+Ugid7sDQnbAMdWH53jtONNLfPK0AWKkzvsNx04ZbCEJ
6orb8L+rKPWA/Bxg1N0X0SfbeEV4WwVNDei1eOs3ILYwXcvhjxOsXkZBIZorCTscSOJZ0aSknJoF
yrpZGQAb+OoiOnNiV65Sf4S4TdHEGGATCFCIix5OtwlLa7X5LMuPJSE8OsFnhjsApfbxPtBQNN3i
RjdMG7lXlNV8GJ/doOMy4r2QC1EHq5NMiNDrHfKoQwXv2MurYXu963EA2ifqkf3CcnLxIBelmTE+
oeUpc83k9RZlXoeTtf38AlnW+Mj9U64T6/r8elIz2B1BhwD/3LUpIUFMMNpICwVt8FlgVI7XSLSq
Pn4dRK8/1+qw7R9pcbT+frYHnuJlIWbQC6SH33iTl7eBBodfNLXAQ5IYo8x39InzX4PolthQhtGy
NJvdeWMCznVvL3wspcS2ajZC0wi7+112yxBbQzYlOEnucxQ+ZEeLXlm3gRS63JHWFdZo3mXtElCq
yfLB8GFZM8VSOpFOdTiUuUi9q3Y6lr9gKLswTTvc/p19gq9c6zMpISUR9DzKs08nMy+yrusfiGNg
sbV61byX3h/OQ5FxYhje9lYlYVAdmsCK6bZiuTB0X0g61cTRZGW+/YaHKXqBRsVAAA1YFhPyGnBN
F0QRZkazLTYo2XsxOkCB3+x2Z6c+ysp5FRCxA9807sJF5ziha82M72m6CtIp+NbBoxhWbsgshpEP
5/fpvAP6X22wJQyeMog1gSnfT7yb8pRXLLZVBlkci+SVoymbr7cH0BBkKlkcb+Tu9xWXJX8ASZdN
NwDh4Yu5Q7rnAe7+b/UHydyqcOND18w0Hhxx8zzyAAvxs6DekGE5DUnpaWZqaGpEJFMu+Bnm60uL
4FUCbdC5VS5Tk1P2K81iNlYWvfnYsdFkYCtN7gVeJLvcosNkm7On+Qq7DHUhi8lOz2g65FwGXMAs
ZdUxtmNdcMz8LD+FtLWajMPDmwqTVJBB8P2X7Xh5Uzltd5VFOdLm1dyQ4PGGdUvnDICybR/OCixp
u62uEWoi2an1dXQ/XFoImz5OVDqGs+1WBY/R+DmYbrPIzFLqtEr3JvcmGTpdXEJxbcRqzWLiIe0Q
B70X8nObutZ0JvBuj7uutvhMpBIiPgxVaiglsVTUUW+IevvHhoTxC+JOrtMoXoAGmIzmfZ3pAwLb
8LVjmP4yF4Ok6vjJvjECUXFdew1xWebVTi3T8s/J8JrvLZNrq6u0yBSveAVGpHNbeu/vqHvJvtuZ
qBjqwufR8dPCu3+T6K1jepIcINOtKjrDIr27MY+l+LEqdYnGYYPGw/W3kMPcdBBZZ35GdrSkae2A
PMrUzw4l5PIXbMT356yRo/Czh5ChawtpM9fUHn/27RoGr3NMA1qRoTaQS966CaN4ZhsewwxjpTL5
oHs9Iwf2jk/N49+VOXLhbLFcZL0PGtHqqnlu/RKefc8IH91QdV5r71VSjbbkX7PKNKIYc3Rfglne
1nm8WG8nN2B5b11Kse/DYIqvdEXjjKnC7t2dg2FXkOuYDToHxgycKVEIrDsgZ3lICpK5clGWaVp4
SeXSIBqkfp9uXVs07lJ8IXV1DqsTZ2mLKKLl3m9C4Kq2bsqVSUgDt1QCpp+iYIHqPCwFnIgtgVWD
5f0fHF4PS4yBSWV56t41iJYxL4P4CgUz33Pq60fF95DnA9zKPrsARblIyPInd1UHanmdf3ljCppH
5yies6KDbWEVJMSS3EdMmQqBvMn62eaLg6HTSIS+cVshRolANEQNQHGoTtXcdps8YEgHUTHK0RkX
Q4/Uzb55Zvr325pUGMjaWN6S9lh0zGqq3tGM0tRUNcTUzkSaqREXC4ApJBqvIGpIsTiwz1GUEAYl
11f09rHaF/ixxDHXTBFXR1JzllYPFA4jdwMed5TLkhk327n/113QDKUhPo/UDkyPEhMQI9UX5S/C
Svs/Fs/SHwwqthvMP3F3aG0Y4MJjUxDrlWzA62o7zh0W2KE95gTGGpvevHK2pVWBb+BQZaNTsODG
m5f1cNpaIlnDRAlKUVEF1m9Cy8XMnTCaqpZLpKTRYaeg4V8/afwCFjEaU1CiI3xPuza1PCwIiGnR
ZhS2jcsQjET6jExeVFOcR937pPLM+VL/vYlk/nSjCzFDM8KW5V8PYJrd6wKlHk1IGC0sijJzYtRp
JmP4s2dD6zGtE130xUHHrqy7lXcGpQI0j7VLwIG4d0pw4ik8JB4EbGatfNW7iS7+M/REUHHQCQp6
dwWCwEv2W9kL4gQLTvbWgm4i2xHsie/ndEylx728FF+xCZivTjFf6y1O3pMreeWea1IomwCEF6Mi
uopM3sJeTTA8TNzxwv3G0Q9dQ2zjspUA6w6iYIEptFya48jMZhnIB7zaFLfzJkMKV4+G/yPXWyRO
wBGuOXri2AFqkJPORwueIUDYnDBW7w+DQAp9p2NxfvK3CZvDalpdZz9n6ZWym18mkqKIAGTxbaoq
0PPy2bVawqLSMO3f4gSfkgmYbPIAB8cfeCpKpHqmKY0TF9qwjbgkplKOLwNnQpf5tTCmMSs7U23E
pU+5uJw5LWYS34BcxYvAhoMoGvYj71h5EVXSULLWV/4C5aIbYwf0yrgJuUBPBGh0IjWlhmT9Yp5k
16eIsabpppnV5tyjd0yqX2ZnjE8WzpTYWxAmqtZ69rU+B2tJqorzffTm0PD38Ps2fbtM74VZNLOC
CFsq03aW//JOxwti0PpSLF1+7MBdYZhI974SHZ2Q79jJeBsP2yxiKHFUF+Myr0HhEAlxWnU/z97H
vwbfYAHjrn9bUrVasQrhAAK7DovrObAXgTDNQLJOiK+h8wMZnUdhJ7xd6JC0b3J+WM+GC4wTMYRt
UNkz22pMncW9N1m/dskjl18s45L7bvR/yP+5kMsu0AcWwqdA2zPT3rYjW7aJkoG43ctNPdRaDatE
jnwbDvO/bsdDr+VqNDEzp2mKzQPZnUqqQGVRCoSgQm7pm+K8+pXt3OeDtAuPQJj5Oou4R72N2I29
bJPNf12/ZW9bsNryvOFlcCzVkTXdvHcsY+/sMGQYMV3rx84ErUT6zX1z7zZQFNTYlck1wtxgxsLr
dFqMJHWvqcsy0vwSwA2DT1XVjUfphxMsHUBf8dOczLufCvNnLrc0x0E1GVO2Ttxfug7Gzc1jlGAg
0dvLc/uFqSSZLGaMbfhwNsXNEWhdQT9zGi8CE4/+yzpop0VolXhGoRuNYtqOLo8yoTXAE5G37zlx
IOjU/FIEr7HOc5XWFwl9+Hoe0Y6CkGZ6vxp0yRqRqN9w3l8jx0/9i0PcjOiOaG0vv4RpEsAP2voL
YLZKtb5cIvCZOcSJNYOK7dCj04k1gbnp9KWN7wT/jywmTqorvREc3EweYm6rXd5XbMXbmXykH42o
xnN5Y/mr8MAH30MJas599qUTxq/ziWVXQaIO1XExu2maOCB8scs1lUEOi8Gapf1CKOXocxIaQptW
QlkXTicQOIkY04JnhGbug10Otyn/NyqZe+HLnTZveE6DCtE5zSsCsSVSGgNKL8w848xHPun7yb7i
n9kvdJdo6qPUJRX8YlIP6eoJ3P7c2L+lY0kTgDJAM1WmYxl8iRu8F9PQKnJIMhdVblidCFClYE2m
VCUckq2K4R9hKhF7nDE33VroBQAK75lo3c98JWK/ykvjjO0MXlNTduKSZj/tEcOiRGX6ujGqDWhQ
VS8Qtrf4bP1C8lTV9IUsUL4qCdnTP3p7VO8WzZ4NK2V6PLIEvHrC+Td70QxvJ8uruh+bHTregisr
bGKMfVJLrvfG91egJ34+EkOv70APsmGJrPCPM1QFcXbg6jHHn34iUwkSJV5IxTMOes44taY49eG9
tw3dGVG6qeN08ixwEv1QTz46QNWF3A2t+6VvPwyEYkSlY9ymUSZMYa/XYTeuPmGc79ToivLxuxN9
UN16BsW5ta7e2eZ2av2/TJKDcs9Zoe6BrWEPOpqtIqlBxQ6xIOeikKM3pSvzFs+8GuDvSLvSup6V
3bmSF9wBhMgQ7MUvhbTK3SkvC0IbzFFEBLdAo9eGzQaOx9dO0rqDf6hNlKLcpArMEfM5BJB3XRUe
F5Pj5Dki/j+Az/DG8feFbJB5Wh3eQESys8wop+TA12bPbI9qMvjzkREQu4eyd/TznXEZJxjTfu96
avE4j/VDhceJwLS1T6XAh6v6KJerY8aeiLYXLaBHsSZEjeAQZjd0B29vQRuxFirGnbvjjL2XH9Ln
5w9e5Y4DvPbJoKYAxjykpJMUPEa9dNd4jTKzzfdSVx+0lXKtGNxPxxKz5G5TV7qOlmmqif44UMv4
HO+SnSrhuVcmYFgkqkZWPFI98HAuexArjgIN+KdOW8/Vwa0WjN0zrGtDdKBlCF7d/pxLnoaJnW7g
r67HlnK6+RQB+omg9XrBMspYC/O3KSGVNVzQ858mcwNsxVZJ+VrXY8U7qcV2cNsawJGjN0af9CCk
2HikhizWAwnt7FI6FbhO3LnkVcHigR87sgFSm3GCNAF0MTVIEIUwSNRraeRd4STcIQM3Xo9p9pho
uBAR+54gqGPopj2r7AN6J4v5jRfZh2Mbs+6243jk7j09a+U7pnKEXuw3oTOCBwq8kp4AKpA+XUr8
9B6bXKh++0V/DMHJH3l+MZdmAeBmM1L4YvhCQbnr4BFbBduQxcvZKCqnQK+rp8I3m/YgYokfn2cv
ooXbc5r/gWOhzjBwF7uUb6T61lh3aHWOHVJm0+dY/QzaW3rZaMkhAwXhJxyqCsZSFT1XWYeil0RF
SBQgCxAJHb6zO8GRKB30ALrBjkWMX2fTweYNjzCpzLPowchzVMSazU4NgxK4CZRq+nuoqm0MAkzZ
0DMCUI0V8XlZG6h5vUxJ4onehTbZG2/fvrBW9nAJ+a4UUeHQ2zbWCLIYU03eSthL5zEJrh82ov81
ujJRQK0+kl1UByQ2/HeKRmmTSezgOtRiSao67NN7uve+Vh5/hHmgLMqARJNPgimDfS4q9uBRk42d
kB5FeBCjXr9QjpjTQtoQF8ApvZGkKZqyMEHsiMwICTYq4aV9IJPtu8YKljbIk3ZZ441DAnyZofqN
Q2PKR1KY9hNDV7fuNgl8/wJvnRaNXdSRookRGlZiCjyf3aeMS5i0dol/YZrYxpiq9tucmy50sBYZ
sSQvXziI3ynt0PQSpcpABTYPejnna2hCwMhOU9puLdri354QToHW8LCm8oZTgIG8mnD/4ZX0mree
rKjHqiVPzQdF9aH3A/31Eoru3IHeGoWF99Jf2k8YmQGfbEukshiz+9dPN9KDP2VZLmJWQTOVM+41
SPfUZL2v1RVDvcMyQBHJwkKfq5c+OmzwlY2hV61BF5jwIuGFVtdiTes+h59pR2mpt1iOSnaeJLLy
hz27RuRzLqsUXyrwc3GnVK1zZVb35oUWWt7kBXCNKKKhDWKhi5z20JjCyjI+ab17ttZ86n9T45mM
b7CUNu9RjOojt5DS2TfveovT7/soP67fnHdFDpf5L+gR3jg/60E/FHvr6pQSsrk1Lj5F1U4fr2O+
aRSLVarmP7bmwSqxm4LVO8NMjKotvpnxb3US530GOuqXoEMr0KGOKim2cR1m/WajwwD0QgypDN/x
dQVW7Ll9hHKnPXqnv0oyOtjcj7DeJriGCkZBahFGYWwLhyDtkuercXHnrIFbeZN4aOSUyuOryhMW
FTSXieBSwqLHZ6HBvRGexUxsF6S8rYQqSTF8n+d/ns1NPB7DUjVzmPjFf71i3Deru6P73iZ/F1pF
vHH1Y9CCUOSxWLWigW575Ph/a9zE/80wXqcIQvmJrI8Y8PpIckhwvwm5Rqw8044FuaN3Imrm/neW
Cy73yPPaZpsO6kbhyFwQ5i987bZbA8Nw167pMLgyHen5U9syzDmz1Ql1MsfWk8TWvx4IfZb3j22m
hHMtD7eZ8K03hkPxNIVUBezB+AuMnW0uK4/VRo7zsL1pvl10F7UyElNT1msrGhxqj0iBTnWj/Dd1
wCuqKTIesi0tZaMqVxanz0hCvOC9xXjyHf/HxMVoTncxi5RCJkZh00CYT33Q/DBEewFGDjNT+9aD
rgDuMdT3ivxTHY6sEQmmkYgI9Sy5EmUWkYXH7yA3XhTgYOwJNkQBbsGT6v4gak01fIW+HuR1KuYI
wnAYjUuNeuN3dq1I37bjBQ22LfZ9RHX5Wj+iIclp2TyDqYr9ExXFu9NPitFue5KjaBGHPzSvg42o
N1MWdFS+qwmPkjVNsuV7oq85XGkqTHB7KNJ2bygMz7IJPzIN/46v4OG3Yw2DVBN6UP8csaRw3SpF
6EsS8uClXYjjly++wRUcR5flgVxMlZhFdjZoqmMl/lqtgSTFd/sv2LMgXj6ku6U3OaNYxzoisYZR
XR75fi9SC6P9O2IdqNF50Kivrnpo8r2x7v3C+e3qDLwLNUS8ZrIMFuypy8zd2p0blVls96NW+09/
WGnGi1fYnAD79sut4BPexoh6NOOcjPoG8qqfnsBgcEobg7TNYQpqqT9HT/mjfzbxfgab0pDSimS3
vMfXiDSQRWFnMxL3tg/YPE96+aaD3LsP3wFhxXB2DCFIZ198ElZf89GTJBNHHLDr/pwDMUZxo7Or
qk9QPRy38SwymVZzn75LUoRhJb5LQBRaxmrSKy8br52ZacMm/MxUzEls/kXHpFb6DhOrhM1E1Fnf
XAEdUermbpKcRRjjucgC7/BsdV1tClNkDjmVxd11UqmZzBmY2JaCpFEluLa0+m90LhYGIJ/SAijL
ZE75tcKXtaiclri1JWsvJ9uO+8/A+gD7XNW8NxiI0NlG7Zez7HP48C0HFtufS2FRuGGtgNlBWi++
Pj8TlXjFAgtN8Q80YzT9gH8u7zLw65ulvzKkkPkI6AkZAuhpyzhdpVhF84p8N+LnNa/AWnJ/91ol
fBkDMczM3x7EmU62Q1vcS/VWj9ylRMdjTUbTN85macldBo0dRjg1ib7im8HjI7iIswuQxs4g2QmG
TarUpZP7kIeYjnHoCNmhvfmXjnc/nU8Rlgn1crtSF+IVWcT7QnlkkJALOMy8zCcUPHz3EYKGLwZn
e6sKC9QE98sR7AD13Wr0Lfsih0PriAd4sGHv3/5OYOF+qC0NxI7zyAEB4opQXzmg5UuTb+C5M51/
hF1SE4Ck0JugxD06j2dNBUfkbCT83qy4DQEJx97tcUqmM41NiDx8eKnp2fwes5QX3PJy3yQq7dfH
DuhV+qXHQa4PNo2lBxMAZTriY0BJXKpPgHCR90WPQINlZoIjnQGszvvw6NMyu8k4uYldxmbdWhrw
xmeDsdcq5MgecoGSSVucX/yPvNPjx1rGVNNzX9v09aK8arHlS+bDosdt6PVu8HEcGVvvbkHQ6qJu
KUcX8lTlBWLDSq7OVOXgv8ARlA7sFkcQglZz4QHHunUM9RZLWlyDlYTa1kszZLn4h2fPcbcmzxLM
cHVpDVjX0ICXlSSrG7wHP7EHRnXp+8rRhWW0M3rmRskhYtA8L3GJrEkBFoct0O9pTtRwYApaEGty
q6CeaoSZifiPcZg0RMYqJ9KhdgdNh0wjjPJ9qutkysaNoqp7vrL+2lT4xpJbVkgAsCKIME2bLLs+
2p1ENCkhodj0bsJNTRi+DyvLchyINho20dNyRSpPsVYncEikpPYzy1es2X6D9k7q8JUwWqpRsDcH
FG+mqS3LEVlAj3gQcc63gF4JagEZt+XLYGUR530EXSG2pAuzMhNWyFQ3edbIyIUQk+/LD1sLYVTt
sSYg7USJ/ft8/2IHUBkimqZVSZdrDLjSxjrTDodWjNXRj7RtG0Knw7uGmaTxWBy+2GLRuTN9acmS
7ZXJFsGMcjmx4BFEp7ewdLPXaYjhwh5mud7W/dS4eMQ2GKAQ3erGUpLkNtpoS4lKyXW8nMsAJQeb
XvzXFgZst+IZF7vXL5RMWbQtiO9n5YvuLRD1zzruxnq0wMZMYHulfEYfdOT05yqx1gInqgdkh0+I
GG3+TDrecx514xZQnRKyUJWHJBMAKD/TCgidKFWTRseGUtu0Z4uKdygtXK/Hrt8UE9RQi/oUm08+
edjjqrE/G/Y/Ms8jl1Q5tOfIYJSzsJtN7IxDmztOKRF28Hq0MUb5tsqW1JBBktmndwd5yPLy2GeE
Tk0Ypr5YbksQuHZMUAJlj+hUpRTbVUkgW9LH+N5icYeScd+y+miQDH/u0HvKn7BoPl4DTpdHFsBi
rl3UO0Z1rKhvHW0c28l8ZJDTqL3ZSCYivGkaOGkfuc+WNjegXE5Sd2aF6lZ9GDZoCsGLVZqPM0jQ
JDZI+hMHW74Q+CwrHdVGpu9hMPG7yyNNnCyxxlyiOCuS/pjv5INWv1Dd60vuQ6t5xh7JaDLayGwl
hCrT+u/vyg0iQ/hk5D2VbiaJMrAbOYsCx4CUfrQqXmO/N7yT3EZqTzcOE2kg8Et4NvBZVZSEoOPZ
XSGPDMvuo0cebrRy9ErDDqXJdPZZBSiI9ssl1xssa104ynTerISREHw7Ph4wDw8VegVn/Kb3koOl
+/s/YwQYPYdMcWe6Ja66js4fsWlVaLmqkqpxrd/JR0bIoW8zMW2PNngKGJS63RxvGauipLfyJRZs
zTT73OBPF14Q4D98VcNcFZAf9lYXdaHpa2gfR8g9av+sQ+Bo+ez5k+UYCuodggCz0K0hIvVObeog
idBfgPwKyqtvZy7+XwI4Bz7UiJCE6hT2nE41lbpvHzYGmP75waA7ogNTswkaek0AEyHtR6VI1Usx
6v+AY+ViKDjZV1fW0qlmglknblo0iBe1QWTOn7cDQ3YwLSF4i6WudrmwCiB0so6z3Ia7WJ5pFyvk
wfFUIjeTHPrvTivNadhbVdu+LyfTaffpe5r//AsIlBJCJDSUFvR9KXV0QPuS9AjLHpXuKmgEGJm/
6q46qBClvAO0EEej+B2K0gdmGF67q8crwtQcdC8KNK5eehyU0BA1NN/n2ygzSdACFntaeR5GaaUH
DOw1K6he6Weib6gMhKBH8+g+aXk+usQfTbpy/mMUT8ddfJnUsJ7TLfj16SMG4RXJE8trtAEb7Ihb
xmhynOI8pP/XAcJFIMSthsZllxq55G2z9g5EXAy24RzCRG2HrqkxZc+klFGlQeMhgDKq5vJG7KbP
PJv9pKKjxZLwHPxcQkmcZG6dVe2ahJUKwKYV6c9clT5QQr/gZqrEm9P9pU57Cp6+Rknzr0PzKZ26
dIWZby/uG330QhCimzopjHhGyMZKyOlOuNJu8aRN5mu5aUK0NIDBasL82HhtbGts+nXZgqrR/E+w
D0ilgRtUKMmF9mcwrrBadLHNq5lYgvFA7G63KA2B/x9qnqCCeRr0KabGSXzQWQfrHzDtwZ87gIZo
xbu3mJVM3xrO/5h3V2DoXBzq/wSrfTkLL90S230MMmSXefOLk0LgdYtzcB+lqKGvWOu3teAHxZZh
lI6gRonaIT9l2fkTWJDIMvAK6ALNiQRvM8LGIZR6NERVxXugQ9O/NXVjyyuYMavAg1S+RYZhbOdV
srpguNIV47u57KPnfFU50jhiZM0vr9hVjIFo0PtXsk4vAlccRHcEMkEvrrFPaOfFt2gdI029ZFkS
znXVOJohhYf4E0bl949LGC/7gIDPsrUoKVmpGdJIe+EdLshLUnvQg0cndc3dv20AtchP4jED5XVA
+kZCeJhhWY/fhOUK6a8ee8+1zO5TjrKmxTy83730dQLOe2s55dPCNJ5xizVpM3aRqH6l6SNkg834
xZsvVcNWRBAV99aDZtkm/wYYq+I+UA3/5+FkDhlJsqsGjP7P0hX7WwIL2zBdEFSE2BHHjnlAdw1e
9iigmdgEdg/3V2RVKg6sSG/eI1QrRLQTmIc6bR2Eheb63JtB9xQMi2IpiCaxNCXQhD//8fZLC4cf
v7VdCsnBPOzVkt+i8QZSI6x3s+/cUyETRSN9FUBl5morKWwo74ldAuKMOXsavAumXpte23lYC5Z8
UGqV7M9jyxMiQlpIHmPFtNJpIR7z6PMFir5XbTPv9+ppmdnJh24bUIhv/LxImbDzXZuuDElyCjDV
CCXKylg5y47LKLDVxyVUurLesfq82gQoJ6sc/BNPbtjHvww8M1Uks+LV+dL6AcoiJQ840M2/3n8i
2UkOk2ohsrJAdQR9pRH0/LDkoLlnpERt4jN1a8RUIYCtLw1oUXo/IoM+uKkRg6Gcz4uXsX/MZVUg
Q2i0Qad66usZPJEiTcXUII/caA7iwxJ2rwHqJXHAxEChaTk4yyzObOE7xXICwvYSMYy+vWlEnr7D
tOED6FziZ5vIoz/nqkod4rGUBHjmvYx8olIqaBGRUzVbaR1RyCf60xUR03qn6QZNzQDLu0TlV30z
2giDV45DSSb/uvj31jn3o9ZP9ggugn6UIb9S3EnRvN0mxHGhcVx5ksfLmGxWmQdljgEX1BHyaSPZ
YGiAJe1lv3MG3fCeoCVJsWXb6O0ID4LZy9O1muB8oIXsP7YVY9o1ItOl2kp87HdxeAT9ptQEutpp
PcCChDv1rqSDOb3PcYQ5jhW73oFtkEy0OsxaoTw1FrMZKWqriDxXl17Cw31mziDaHpnh+oOq0+Yk
3GB7V82jTesD3JqHmAsQQlB3UcK58YnL+fPTaT3+V1GTkThsTN0dKc4Ho4ayZUhhIcEisR0rZIvn
ucpD3oEmrCOdyplTA9u7ZoWj7wzm0iPRcinBihzajVCuJnb8AJL1jev3sk8fbiMaJ3BzkK4KnRL9
9eJPboSq05cqbB3sGQJrVDXEzymYSJ8jZgCfpz3KtG6P/B2UTvDJa+/abICff2BG44o6NFaMyWv7
7m1C+unIB9IlS0mTdjGWE4WivMhQFOM4s1/Y471ejDu+JYlynYxKWiadPQWg9wUYhLYahh67ksDQ
xrJ2v0JNjWiELOXAWP3gvyFp9sRHVYbu/gJNqN0wZvr8CxHrsnHjJT4nv7GMqSfcT9SVaDnVUTqW
kldSU+H3k9GJs6ZwGLgfbhP/hbdU1gZXbqPZWoueuthafym3KU5obYk6iZMjHEfQednmu+0YZOIS
bQ/POHKx8Wi4ZZfV7Y07dCtfLVPVcq07O95meob8+dGJcAYisxmW1Fctt02ClczIzmwavYKD5816
oAsqrDcKQLdr4CCumWxPlrJVJX4EEy+PYbJhD08E+8udgFfNoJWdxDtguE0rCShovmgKb+8W/K70
ozfFopiUG6S/1GMmHYQiiWAHvhU1Ro5Hjt4qNxKubzXznys4okTw+X+IBMeHwFDR1v5Ub6yZwUWr
Qvg+2pcAUjJP3bBKkOZYCf1c4w7ob/0z1ZKeCyT3sCTsBwu5LufUA+CPWfso78+2cxDUxzpLWO6R
ZP/1iWYwxR43KxTBldoaAQTTQ2iXBNCQsJ1vTPWoQubBt2Lv6/p6NFagiDR8S0Vaq9zdCn0N5GTc
jpZZXR01SQaIGiwrtcm7uwucwvuyOIXSucz90ns4ra0mJ/UNq63b5ZoXrioNvgc1Y5JBlYWNLQ8q
QiwvfkWTrkhvNe60yYbTFZmdMtXaHFPUG3+jpM9Tlmbo3IRz3CZRD4DJq+fsiDOC8ZZTnqIHcdZw
bN2XT2tkM7coXd1O/hiKVFK8JRG/A+5ouDCAg/u5vPpkMJJ7JtzfE1wFZZTKWjQ7raJYCwWyytwz
vJRVkhZzl2qSdKuP2/EPOkFDlsX0lvsG7bSbkVdJAUEZz06doKqME6xnm4HtdCkckl5pwNIlHQd5
kyz3ZxVof0euqfEdFNmDjtKcnt5YDgubNKBDSqQKRzSBmwtw8Di0cwKTdY6yd+TLMBTg/WrgZfWA
aB21cexuZzyEOGGiUx+gfQ1nbAgzc4kFZt/l1XRiKUuUGqGhjEX/xrlvmv/ZB9Th4bGVvK9HTqEG
zuXkw43d4i9tNhTEOMDeFmY77MsE/yuWKaF4kgL3Zfj/g18OeBLPuvw9AmrYXOcbaDyYo8WPErIO
v9Do6rQm/5YfMvzll9fnQsMJ+CnYWzJsd1NqIXJkKbj/4PgANRTyaWJoBRfgg0jLzLzLz8Mh3zyu
i6yjZ/FiiqKpDCOydH9ReOlcnCnkttypCnA6cVJh4QIIFB9h+fb3rKUsjz8vbYvmgwzNlRfaST5i
E++KUkY6JIQKcJZEqRxVc15evbPvAG137U/StqY2mbIxFLIW26LzHHCXxpm2U846sMRTIBjwuBoh
yTOcxVvOyfTsKdJtUzKIi0qMCM8LW0wj0xxHmM5Tpq/SIUUxIlS1XhziZfomCvuClIBK/5x+8I8Y
rDaIWtaKbzKZuAjCoa9c+J+foq/X5B1HZO3wyTo7OYB6QO8pDZCbF+h33I/qdULsFh7LrBNJybpx
RczNVxPrAwDRuduxW+YTSnM3KbZI75/GqDHos/Ftx00CmBF9Z+LTXUz30UGNA04mNsfOtperQnbD
Oy3wj5DsUmn66udpD7JynHjI+6sXeWokPXYS7lhs3SmAXwyGDC6VwnjokcbyaQP5ow5Ed5q9mkuM
CwoPwLeL4OF3SqlLV5x7cCwRGxtsnrkWW6SQiLXb7bzafQwx1ZICZm+XGEupSCZbDv6cQT0gbdoy
Wav4Ezt7ZAzA+wMlflppAfYm1MVNqbHmjRf2mij1NdsZXtoYoPNw2lue9dWiqspX8fn8KeNQ/uhe
p7C99J3af9M2zzKoHkXmICA5PDzaGsOGUKu4OSixAz49PXuVOYtEAARW4wNQwbgY5mCeP80UCgBA
MtXZz4PZ9VbHoksW//hAZnpsSdsc8TwlDLNmRJZeosLF5AW0+hnLroPNpzB97Pj2il1fKsBLv9Oy
SEI2gHZrEz9Mfh3avGvJFonRbRu5uLSj/48DzC6dHIHGFap8RJxHWEFFE+XHCjDsS2ZCMyFUUHH5
Km2plcKj+aJ2QZmv6FC8PSYIOjJ3Yy/DX7l4PfALr1J95uzqce4ju2Beoz/k4vmTI3oKZLZrI5mK
a4aSGM1PbTXXbjwUFOLxsHWHb5rZlM2uuc5Si/WYZ4liocRAxnuWk5YlIiu5A6knaZhLyI7jre8P
xGHL4trZGgzQsuEUErMHTZP5wkwAeG4Xjs0u4g2RBkBZJ5iTdMO+rhgW7g0kWgXZ5II9NCRo6BD/
gZDPc65qibv72aOYM+NK7z7S3m6uOPyxj2bt4lh+wSijZQyjsRlHKQhH8hh4zhiWgk83UdwTBP9i
1UAJHu2j983E+rhqNOvL3pR/O28LIdfABNmcQlUAQzbkyh0ebg+qkzNvbHEVSDrbyn7W+fKFtjq1
i/i+PVAbc5cOksdDASDaPidHCgRCooi7/0kcF/CxUKq0+7fQU1LbURACmBXT3e3sWA3oUnG36yg/
oNFsSuS8Y149PjnwlC7KWSlmK8rmrYNc1J4LVlppd5hfMEOdbdt6eVHuBuyH12pvhxqQXCLC6+Ix
QDTakOpHJ5hX8CYrvOdMc5ITXhWtVr/HqFBt8m+8SsbxsPT0IjFRXx2JEeKpPR9EDVLLa+D7jKiG
PA0UgO0CEDVciyCay/QvxUE8/VC0u8M8Y9yk97B7m63OB1AMo2z2U3/lr4WoUXc+WP4YCLM26xy6
hDpqBbWYEaengxgtbHQW1aQz3N8lthn8SWX4Nxn+g9Pogt5P8COpxm8hamrv9ywqfQvezzkEx5sQ
RPJ0Xo9pJfWYHSI93Dfb3xQVr5gSA9PSXHGears9MXFX7ffAZmp5Wf5w0KJwfefyDo6uBqcmr7wT
MPec4hvU9lYeLYpQjb0qmO1k+ZCvpBc/TOFd+4Vzg/qs90sGSw2YOdBPGyk84uDiFH9JVLv4+5xZ
uT+ca4aPU6kiZkadwsLy6CnVQ36LBMM4WykPM7SlV/a2O/y6kkGcMIlr977R7MDku47X0DWE93iA
yQVAjZY9FVPFhwwBTioo5B2yyScAV0qUWZ9GGXyDBID6E4DtwtGyT1zI44GzY5q2rVRQAkdz5b+8
+JQlgxj7XQxJ3vnYwvox2zIRQa0mG82mkZM2ghve7T+59fodRb8o4PGUuAl51889AHXI8lj+40Id
TeBx1jW1PETGkBHnzvR1Uq0uA5EhwdBgknVVFWX2C5kFUh33mi+XP/YM9nMQvErcD5I1yjwiQjx3
0sF3gWtsHhjTH8u0lo8Rq15d7kQ1kFig2ulV5cW43PEJLsJ7FTdFG0yZ7V2ZOzCnqIXgYITEw0ip
toFq7jEP5FkNaa8FtxJ6XAROTsME65xv2wvaICsqO2yckmX34Da3wnzWdHolG+KvciPiXtjdVjAV
d4waG1krqJRuRSGahyVw8Wj/HeKlT39xWLRyMKVPJ8g5YfFHq+NZydrABjwOv11PvrIOvDpN0El3
pqwf/+MxZfQNVPES2VYG89r7UB5vp65nJacnRntedKF0OgooXcxbwQH/HYaFAAAeftK/rRkASMZu
lPmoosJ6l1JmjDgun9PwxHJK5rXNFpA8Hjur+7MKKuD+3fSPd33OhZ/HRv19JF3qTgT9bvXFxR31
Y9j2SVvmzdhJ6XQlZGW6IzYR/kEUV4rRXQ6jywahrlCm2c36+Sc0JZ8+4hyiCPAmUpuL33XO84mJ
R8imntaWe9JsA5t9qcbIv5SgXWwXo3gnuVApP9vGKINwcllDcasOL8Jl6L2XqpaEb7dJrUZV3c9S
fGMKn33SCs4/u8NPjs+K2dwa+u23DnFgKXT0fXtna+rT4yinoc4bhZ2d/N19smUqkDmFNiznbyVu
EleYNfGjkN/uuO5UAerb4hUxApCQ0yktR38CKDeNyrbZ3txnkSvpEB3HDFMCjxjVbkEQfSPQTfoR
WhbHk1bxkQiXzX3zbZdZXaZ+ONpqQ6KYRLMuVGHbBrSG/GGb23FCzOYijqxvf2q6V++jyv1DxaV3
4he9ueFFlhZa9wlqJo2BWnzUsKAyKBSGtl0dRFfKbAreDZiFGOwOIJXrYiLTgWLbo05sP3VMv5yE
YVQFT9LOg8aLydPToNsKG3bA37hpCufiThWfP3TAawc/Nwfjc4Fls/xZZHt0WrNINhR43amne3mO
Zo9jpeq3vHaWWd5n/W7dEDHzUbjrV1oUoWYvOH1Wp3Mry+ihPrZdwsIqkIJHqq2m4RE+w3yeMoDW
MGFz7+gXkFwF/QHkxtoMwJP2E+sHuq8DS9R9SdDB0uP64hXLee0l+lB4CAbOHlbhazRtjwGqDq7b
22PsNAFrryQS6fCXRFH5MCgAkp1FQ0btn3TGnPv690p5UnXQIpVGQK+b0VC/B3yoHdyeH3vnM9Ej
R63u+p83zVitDCEFukGqigz5DXCtSRSPrmsCLka3CVH7it2FbmZLMm4MlnThWy4aqVlr9l+RHTSZ
dKyedUjKcY6J+LnoFiILKiVX6KdoSLTD3tOCzAcdtwGPM+eDf3uZR3K93eXVEoUMEec/OgXQCi0T
hHYC122jgNKJN2JghTCu28iyNHH2s4tpONMrAEHsitCTki5Cb+AwTwiBqpkO1B1gUIyq+ngUSEf9
0lYxy34IJt2gROfRURQxLmmasemujyTosqW3HmB4hxM0ZuDx7PQDmUi4UceKiNqH1eJg8Xw9h5nQ
uoCQF4naCureMHeEIN2HBJY8MNX53c81RqYWkiiF7eq25QLKDbBm4vFLDBFHjg8jFbPEFKvOAlqW
PGiVTlK+8TVj8UwP30E8NamSg2Y1IHoQR6tiSF6pfsyopt8/46Eef/rd2itvo0Q0tGL4mBJJ595r
0+LQ2xSKSGHH0Je0yOQOOKw3ET9T4aIyJEo61CDaFSbsXEEp2Tsoa2la/LVvmm/SQ5Kyzi7V/Qeo
3i3I56stpxjeZsVLptlxIuXDnJ4jFaJn6LF7pTFoeUETj6ELoyDOtHt0fuY0Xv82RDkOCaLQwhS3
EqyDfMpdm1FIfGwtvekPanFUBfcWtESh8IPNVJyG8qOBIXPpGRv1x0+pGyJ7L7SzGsOGlEju6x2f
IvA1AhKys2jTWuSq35BGGQbMxgseq5AU62uoEd8QKTU8VUN+qycgCxcXooWiE2b2kOQniby5h5yQ
p5ytJg129it0tnu7Prw8nzb/YihwUSzy4LKkk6Zp61UBL3pSXQPpOsx1+uYSCzTSdBEszrPmOJYg
/jf6QKzlR6pf4ryrPsfVYom/3yabdORJrIu3hYJfcLVSb5PzG2SVaVd7CNqRTU3q+uYqMFz6U24U
PgvoZRKq9c/yXTd/YEZS+dcjN+7n6ZZXFoz1aLuVSrWoVatKz+QWqI14VYsXUw4xudtuba7kMnni
W7AjCGNd5rUVlOoFuHQmpxu30Q/YWwNRzrDCJ6wMRiSpji2TeXWXLWUqMNpKvdUrbWgbQSXOdjVg
QWW9ICRpraKklDPwZg6MZNP6SW1XEmOC0Qxsa7wr1ntnNLtWdCsJgIiHUtriZVsIfdCGuB/ZYszH
qsFtbvJ3E/AnvSVXL8S8oIznvGv3VFvs6vblIqUxV9XAMs2VVl+65hi5XH8Klr9wfZ+NpWw50QX7
D8zEmOPJxasZ6ZjnoP2dD2QKnZCNcl+vvJPZ0lJTEqLNGSb2Ya2uPNrIEG2/tzRq1bs4zeCmPt19
ht44qR/hK4auTaisi6cNnXCklWA0s7ySXPzZEqgrLinwaWpSl6qRm8CqXz60wxW/T9CjEiEud+rj
poEBRfuwRLrx2XT+A9ot4r3BnzdKl6QvD6ilBGlwKTM37REBfCR4DxJJl50kCc9NQ4Dhg0aOuKDy
1MKdusGbltroG3BAOAlDhRhwkI7lncs6xYuRbgkkynFYC71aZLeC0LL1JSrAu8sQ155EIMZ1XGr5
x7xxDneBq1WYgqQrRTJ1RURS8d7Cj8V2k1cOVS/Kbxxic5Br6QyPNmPaoPf1TH59ShXzc0NawHiW
sHwZAx87E2Ul2XODl9rZZQch664vJPcQTg1YXzVZefMWCGP0zlGCGYKjppGcxB8LxMNIiECLjJt5
/OiMTCOFTw43aYAo9iqVs3cpq0u7QTZWdM97dQAvBXR0X91EQkxIDdVGpRqDPpGSZ66WOrjolVE3
uV/b+Z8Brxyll6RgP1PhsvopC4yTMbeANEa5FlvlAOTGKr+p2rKQxFRWqJWwqDas0g6qRsz28R0D
dxfk1b8L8bgA2DrhevAKDln1mv21e44UEKmN5hvXSbiaJjeYRYg4lIe9q+c2GfygWiaeLW4D5dSl
TqNhGaOJv9h0I26fDzN8Ad3bItSGJTFXQbRCqL0prppOYayMwxr00s8XsfY6XNhEexDPqIzEtm15
4QJiWbXqBV2fADT4gzQp8DGT/P7dlwh3EwWJae8Slcc2tMB+cGdWun8+yx4FGozkCBedHr5NiNar
6hcKO7WSTrHTE+BZFT3x4/Gx1YRAKKeLaARqCXPTAtn3dsTSdY06flq1FhebrdPvnWjKN90fY/uV
EYHmxGkUlN5kqMJzQtoS4fu3C4nZC+MkPkwEu12hOXKdGYcjWyftoNpr1IIGeMUvYKevGBg5gsqg
rsCQ3xrKXh7jXC+ljQzyhCHJnLcOxs9EV+GlJMe7u6sT+fRW5a8E8rUeiy9HwDGT309MWRERgj5y
gJZEmK3Xvjea/IUlyvjIIjBAo3mzGPe4NTt247umwK3RS3T746bOpLNC+3Z052SiH7vUFJONEaSb
+xRVo/m+UyisAJftFr2hJ4Hqo+YezT7o4tlRPtIxOTh1a1iX7urwa+qXWO5AOWnpzLnxy4dQH84L
PMAaciPC1hAwOrZBVQ4s0gKH/1jxO+nM+jM25vDwc1fa5P+M6YwMDtUY5jmHJHf61nwBjTSUM+V8
EAxJQPuxi0odVMy85UgfkOA1UGnYlre+bfMo9qRBzsO70ULVwsjDIwHiGXy/rls+MT2qtwD6zyaF
06991QaXN3tUx8wmafBxfAa8UeZsddbqdZn7wEM4TacNc6vOGFbSf0fOEAoM++6qyi9zpD1fDTCq
ZJVhwU6Y5GtffI9U+/Mxz7XAMmEiYHpDrhVqZ6tcar12y/7cAyX5W04jbuoYTDJ7NnAgFq/Iz2dG
aJRCxauYoSBa/IBWCnfotecTHU7hfuSltm9cjZ19Ic3egU3/PQf2FO87T5r+GaYFmqo8gN/Kw9iv
o0T4TMu/qwB5pyiKuvFckHbt6OBOy+DNXPbj5j1P4WUz4SlD8i1o4XxQcHUqLy5pxcLRJeS64olL
5T6ucbsmzuHVhLwzmySg83NG68ZpWoNbsljn7oBNxdrXViUGBV7Jyv5l06FhSPHbCUvVvMcZyptk
dXchnPF5JWbriO79hCW5gysJ4iXHdf18OnuuKyivE8j1SjEVFrML+hC5qZ08Wx3+gXjlINECLLnP
1fGdmzatGx4pnezjwjhW6hket/Fp7cIZb8cQcVBowF5RUaSX1MTWIE9SY+5CCoQw8+adQAIl+RUq
Qk1hXlbbPa8RjUCx3ZUsN0JQ/r4lx+1fsc0BVz+jGVgUKU+NPM3JVL8WiakqUiiqudlslwLoBTfA
pbuEQifR6dlqi6cMmV3AunlmKxxL/3YzqX3RA1XYMTkwb1hKDJJr6J1UU8YkT3pbXwHcilQLvZyT
XjdDrDAgY4TSBqS8TimlptmaEOY8FVICl3zMmJdaueH1/sEbdc5fHUQyV6BtmBoxaI5MN5jK7L1V
GdMfnM517QHsNxKYDgXgH5vBgYMBGSRBT7P54rV4J+P+qSnnMTTObyx+r4FNROgDqeHkXMyeCEph
X2InoO00Or6VoAePE5Z4h1sAlhc3tyDfjvBEDwCYV60p6Osw1j6nZqburAnFajoAxx14upLa4fsn
PD739jlbh6eIpIIDcRXGji13/+J0vSPNs9jUVlxTomr83o+s8Qjl3w5voIqDM3NI9EwUM2NVFwI7
Rh8pmkNsGuLJN9N9bl9qXfF2HtdUKqgmT8JaXsoBdS19onzE5m/70xgBWzQ2eK3adEFkrFKHc6wt
aONB0vhEPjPQZymk7Qfr7P0aRcnXSDxf7rw3t0CfayU8qVHGYOVQxJ2gOjsIpxoJsfkFni5y804G
lE0MUyh+2LQRoaBAoRrAmnrfIXcU12j3PeDu46dI9+bTzjfoSNQGiK8ZcS6hwv4c3U//BC/8jSmY
BxhaK973MN5Lh/qEEvBtvGYgT548uExY81vrdHmnvUbJ2JRYUGsGZVszxBV1lSVYXCn/RTxt4lMw
zZ4ePYHnGReZbNcSWD9Cdc4+rcuCo7/9J6H4NMLEahaoB78D0ZtqH3mlXCUCAPcgF0dtBmUYN4yo
tTOrttqZ4/Hf8iqHic+N1lZxx5UGmBQ7zGGPPzOnGSdnltWSRGA67sdX1tFYSTW3T+AfpNeG4QUr
Q2UIbeDEUlhNZOTafP2/UjbWQ7VROtAVoulb0EjziDX1EvBVefTUJ6AuX1u6vfejc1OdUioQBMNy
4134NJ+xdYyOrqfrNLApTItcviTnIBnfw4dP/qDOK1pA3heoffcpd5QwWBel6/iZEpTfIxYvbEAs
1+GL7VRmjed6vRQ4e9krknsZSz0SNGze+HAglyaQsx1404yG/xnKIyLzKvg22JFPuH1GMxvsu5Ny
EtjMaJps9xobw0vbxRdGjlVjjtVrK4EWQiEw2zgQH/D7uq3LOaOGLoxCZ43Y7hR7oIN44R5oLYwM
3Kp1f/cEixH5WZgAyU5IzYnMdUN9xap2y+WTyUELTCnZlWhIomFHcjAg2FdmwIaZQrjEKXai44JD
mYsVwtjzznjIvcPToxXEz6mxLjgP8UpjPy4K36+voQg1D6TZw3l8KUt3NZ1uZ7WRCdlfaDKKW+KZ
+dYkFidIxucBzgXWkEx/2/8SFXmbfOzMJfaBoX9voq5KNqL86yh/j+gfrTH0UIlGE7anMg0zDe+h
zrLVD227WjytK2z47kN66HAN3PJwVsocth2KhwiTfAOcROxpBc5y+jxRuotjsfCi5f5XRasHpA2m
3yGRTN9Ax2adTJVhN3dGvD7AlxW805ABtE4jzt+HSCHFFRcB8l+yQgEHtH2Bux2RgL5dCw5N/ztd
d+XFuQGlBgWaY81VxQr/F7t6HvGBVYr3cAQ7lOuITE84iNEbWOQnwTmemuDL/IP+a+veZUVQ0GUe
5iKg/F+VThwdqMSCkdw/fEX+dot2J1VHx032AHrW0Merxy6cYbFlTb2iydRK7J7dhNUZfBEV2dWq
nTD/8fXCXepcIeG3Z2PfOs45ks2xJcF5E6bKUpGfaDuNaut9Tcq8q8rXwDpzBc77PMxEMvElP1nq
gfBfSbitoU47ppAdTx16IebCEk1VqQBcChAOj51gOqPxsudlf+BXwv2OzG1KISXjbHvuwknBwXkr
x+/nFa8q/3o3sG8947upNdKEmygL/evGxO60IPmXAWlKkuLUV5flIkNMz0YhkUuybfWWw16RgxW4
aSna+xeMpccmIoTCghRqC+5jzisX8B76wqEfsJ/bsNadmGiIhqS4Jy2gBa0PWRFJ23tumsXqD8QR
MIBm+wySHxSVaWv+1e0/8f3tqAYtoiL075EDt/3ztIJgC5AGBW4rI5x8yJvllmCM2OdBngkoL6gr
/4xOyW/HFPq3ZtK9a4WjRrSjV+omaRWEKVbwxGeQCBlpz6z/RG4Esx/DSUrRyne3qwfntQa7CTPy
55ktQ3BqKCATi1Lp21cPA9b3JUqCNGHHosbeuDsAK/Irdqkbo0ynpk1gOXUPdH1SslSrqyl2q3kE
kkh3C+cDQlZwQl9iTzXZgtroq33pdiDAxQJfxLdpAK58QdL3wq49JZ+yASkh1liuqXbrK93VJpoz
W+5H8HTPKuuFOqTrEz5LgMn7isC8b1yg7v3Ba9fPhJzZqxnbeQP/Em9omVJkmKyhToc8WmX5lSXF
GYHL2ykHLpxxqR9ICvjHhjGqdxysLtnlEZrdkloqsBKPlIuF1OtCJ1Loe1eE4CTJWkT7bch2zRHk
oQe/KUTM90czNQLkpvVxs1gehwD+YzK1ZhXgCQdmABNU/CB8qG7ChtfexcDoRf4DIMdF17DXUMIi
VjPA9y0jmQ5yuKc8gBs8wU5pKi3jlGeW0TMto5a+GDdZaxMuU6M2SnxYgfysi4YbihunRkZGf3y7
WJib1x6Ko7VSJiPCQAIzEZOC0RQnDztCoICqpUwOVQyi71Ka0RPizxjjpA9sO0JrN7HmKBx9flde
vvj7xJVgWRwB/g9RyT419r2tFFCodaFd5qBIZEmsths3GCdSNbKXqk5qEqtlbX7Hq1fDWaHGXaFA
ZCEPJpodOsfSf/2gf4D41/dE70YVGMKTdILELQs4rvaMR1UCwy7GBMrCyFsmyrLsdW7YuKDDszBY
B7G+QX3X24JihHM3KPSi9z/ammolz8z1DP97Qpl4ljtdG4cpf+FW+txtlBaN5Dz78Jz7+l711YP7
7hf3Cw9s7jUa5iBA7PpelgMZa2AhFOW1dj86wnIhP5IXxSv3OV7paQ/B3JuRb0NkKmlX2UbPIjhz
cSGqKOELUFTPUUB4Qj28zgDmryWB7DuEMi80PA54FRRej5L2mTuUCt/dxIZp16cOPR6mrko/orjb
iYFkOQuEyTGBuA5OXv1xxqsRmESjSQs6fAL/LJAQMxA58NCZZyWKjfOWJNzurfEt0jYB5V7zy48h
OMfbP2jrCvLu2ZjOT0yMOEPCZDLxC4tfis5yhB3EQtTjk5yoDbLc5dONJ1f5LqaVBcB6JqendG5a
3oP3CzMUODzUH9AZwppQyj9kaXUunMjC6pOZ7s0hcMEmSwqrqIHd9nICr4+qB6GQOnPtFswHZnl2
QBnJQmoBGzt0fFEagvvir6ZY8Rii/iWeiNYZLpGUzbeAOixQ/Up0WqPAdnezd8Vljy+SzAMSr1BX
TteSqKnw4IEOaYaufA7/Z+ONQH6n8iXauyD9VLWrNO9dclcXwOgEnR9kXznS8copbuKBMBYm5RB0
nN8G+EKMnBHlq8jPqr595xRsC3KPZwlR8Kc5dp3zAUqA6pC/hmwhd7zqPtsufIBm34WR+I4rzEFD
ovosuOYrpq21OWdtqkp3glWb4tbmMpwck77SIkI9Ue/uWveSyOcXhPD2T0oIeYkkmtXXNyar+EiW
HFNm7Jk6SB8kGtTgnPADb5yWiuNAc6d38cUvTucPYgDSR7QvAKBNlUruMbQbg/j8wXMebk/rwdiI
/3VKqBdSk4SsFtYKC0xqwiJvWR9qpjTjq5Xzj/FAXuZ76JqKFAbKcucz+pWyHN7dg8ntXvKqLqmh
TNRqF0ZnqxCZaj2mALEYc6LNlSRsZYerYaNXNiPiszygLtxS9hKDu21P9TryDom+E2J3G7Pl/oW+
7uZzMLfoujLAQpHZf6RVt4E3Lvo7xcUMeeNIvXQzfm2gCYShxLWW2vignGcfFQzt1vhBkMvrgypD
Cq+7iPuVUh92QvudDrGwdmxVx0JkAV/7US2kRilOBxInx+cGIfpTBQtjcyi54bKx1dZYgjaun1rA
NugL/E1+R0R0N6ho4/pODf8BXnLANeXrI+nclgxQ17cFQ+GHkTmTiqBjnnmXp1Uj8rQpwJuaGrZP
AxZvD6Mka3iCAT1MMrzZ6l2Vqe/Ehsyzfuwh+ZNozmDsAIeSrk7q0xR2F2EYQjG+Xl0N/JtirGQr
QqkywwD4C3dFpo471oYkIdu6E+bCBNJEq2SFNRiAVAERFJV1zScnYWBKXy/LQMkNMRguBcatFfwT
8XUicpRx+2ILZyyy2/b13YVBOVIh7vq2eQjysn0iNxPydLnacGGMCF+BE7itSaKo1kPEN7ywcj/7
9H3QZDLAKcxEJeCJbFpU/J/bHj9pjF/7D9bkcY5igHXULHE3rt/ideMG3l9GHnoEI/ohj6vf1njF
HCBL8LL3vDM74ax/QGH9ASqxduxsVkagxNPFbXNM2Ue64tEYJ86KwmFoX09H4bPJB94ZFRVqUWVr
VpZTFu8VZIlKucHbP8k7c0YWxDPbaVE5aDJiU1AI+Y3i1w+8EWvcUFi6Ko0TLshyLKPPDZq1arT0
p1FhBxGOavBG1aUAIu+3np0QQxOZOMHmi0x7Ry2SMVrQK4ZIxa5mkNYZKnNreJfpe3U9Kj/ZXmR+
tVyXyEDOHWHBqULPj7t3EYb9hEJDvBo7zpzXovDSEyPjiqzWT9Ifupqcrv87HPNybkLLCyFnS1Gr
HRHO/Ms38vkDgXHQ01QeiKhCNuOWApdYhVRF2Z5s8O8lHC9jQuLQWP5/0ZihSB+oa40r6bm+Z3f2
dUySIPFSAMfNhL95EAGCS3a4gtoIBaIuJX4QjyW8aUIbkFOWRy+Fb68y/aU7frhso/XMdGThdUTq
CAt7tNrA688Xu3vOn895tpIU99c34Xr0Ki+PYyoO/1wXMS0vO1p8YxHXzEJqckeluWbNkJ80lUVP
mWQ13zQq5TYmdW7tufdP7LuZEQzl2GQyX3+IWoPklEDZKW1FJa6cZ8Da9lEoDvdJ08HRfhEKZj6C
HyOaOO04dNt39jtugFv/WlvWB1YzO31Mqe4r+OdcBPtz5XBTjxcPtHB3HX6JCnzGmsvl7OS822H+
L9p3cfsfy8qv2kdivKfs4fPD2I39rQXRiyqGIvd7ijaxP3HxkngXmGpINKkEGPbJVwJj2gvUJBvh
VhNB1Z8cFRNXjw/3Chtvcu1AQREwXNgLlCdpNXvDX0NepVl0RaukeJApKpMSfEMStDID/h2dGUyi
yClmr0wMvwGHo1BZ98GF19y4whr6i2GtQ1mH2oRMMpkZgPliTjY/6Lnb2Wolw+xd2pw3fpxhBpI1
JkAdufRVLHQwt7NOIrwEBeeL+7nAP65+j50i222dT/Erki5TEpIbjB60BeoXoQbv+LhL1emLalAQ
Mebq00/AbGwUjA+zoZtLNE94rNXSdllhzsrBV6W9dpxPFiWK23hWtQQwRtKPUBMkwU8eBfvZ/a9M
b97Lk6m/q6PQH09Mdzao9iyLlET1Df7q8kZC+54R9fqPzWIAq6UTcwyYPPMys7Dr9El2FkcapgGw
de5hnSqp5nExbs9WhJZz7X6P1y+ZQwY+vI37e5G1VQ1fQhZG/bPD44JLot7Zt8BLv1FINfZHGzxL
CSXjdJ2iT8doGQgei4eEUIN145QkwUZfB02fOm7A3pDaAiytCP25YLtx7c7dVP8Z+upTRBILEvlJ
VaeUT4n5tt02xpI/rSQ3w58mUDKWVEx+WZQr0jqKv4Q8jFGLmzpQ4dxP/dbiwmCZIa+roTI1A/Kg
0vlfDkmNwk0soQ/q5yW2dcrAju8+tc4uPX9fXxY7cIh1KwiZKvWz7s17DzNmf51bLBxAyFz4bxXe
+fekJCj1ntgFiaIdNcop7XhEh9EtX8wJ0vnRVp00yUx6ZbIwPk7fuOepvVtxtHoT6xO8bcjktQDS
3GQPEhd47RRijImytu1dj+e/K5LcNTTIwaXo3Z9m9HCCMxFy6dPtTAIv7HOc1dyFcsywba2xFf1Q
FI7uOcOS4aBS5vP4XcDMQkrQHH8D76+ImCNLGcDbI/VspSRmq0PeSCSGpsk+hiJyrOa+RfSl/4qH
iaWBFWg5vbXj4OfL00rciUFW4raXn3t5kbgHYUtqw/PY42xnyKEj5/KwrTuXZ6lkM9LcwHp/N3qh
ac3F2iNvLEDG8515IjLOq+tKwBx7d5jTA2TPnnQfGiZoaKK21Lnn9pqZq+9MGzaKtuoV8sweyeS4
K/NwQ7LgyRFG66yEAd+IPiCY6wF1kgl3Oe0quNED2WWDRjNTBn+XYl4QmmM673vsEOKlGnhy1yk/
FdnAggQFqu9vhXSeGabSLKDuQ+NI9ptXX4kOAyg9TqvnIShRo80e1Z8dUTa1mLZw5t9OVPC1nCGY
I6ko1em7k7GLeb8pArSCpDLmOGXlr1X+Y7xFLV13EMgSMrv7gS6U0Gu3RdTbG7JsPfnVnN2Dm6Gf
Dyc6nNtICSKowUmu6QP5h2Kq+7wrk+ZwbQmG1sAKjAS7Zp63NGQ6aVSpljrP/zNCthadrHluCl1P
zvi7BW95+6wKwPqGirPYxs+NHKLi/KGzZL9YPtKrVBLtmCWyuiMA/dBw72x2ZnJLcbtFgCqHOeQC
FCzesRIUJE5ZN+D+xgDA3Yf9L2HrIPvfBFCDJXv8WzHchpClTHP91cryG77qeCJcvrA/L9Y2bL2B
PfNkI845uNGIzRVKjl9oA2C5VUxPkP7z5Ruwuy9KCxkief958TLJLKWmH+IFm/oU7bht85h4iXB2
rNoTrEC7NcDhen03pAxWy0+hIFqMiaO7zZ5Q4snHW6KNFSdXMtZuhdlxmJZ5rhoHeDysKtIIeGRU
iiDkxJrNm0l6PYRncckPFmRHw52X6iWRDKR0+/hxhsGksqr+/G9hlKHDQXs3s7UKpYoFV1zqg/9g
nuyKz83x7vRz0FzOY4pHFRINgxcya+DImU2I0HWdrCgxHD/LISMgJw/OKX0PwYTXvBGUfWOOVmCv
DBCgPMVwgQxfvx0XsaYwSOxLo9UkebETAUPj+q1xDz4K9/jO8w4+l7J4TPZOjYkK+DwIi5YMkFIm
7zmPR7y4jhly2J1rLgspLk2s7IQ6XlLki7LTYmbIbfc9DsBHreISJevdKX/SRQTMoSkDMypTSv1V
mler96KadowGQQ+aqX9JAIJWHGMLXIubabwwq52ouXPLwougjR9bDiKo2ZcUd8dTBmhyV14NUj3K
dL2FoDxY15BY6z/2gHVYtiasZzuLt1fzF7VEQRa88oHQpIbhI/yfxpWZlUogqBNHXSSZ7FjmwTUO
bMobRm80YwypS6bk83amaRw0Kz7eqZc/LJrnRkmwnGHp42HrZ6ua/WJtAknOfNfMWemb4kImcftX
TLoipIzSpUMzove36hkNKz5f7JWVeAKfN1LXhrtA0EF3fJX44mAbjAEQwVPvl5uFEmiI3/SSpW4R
pU37CHSjbGdnM+QL/97UcqlO1bMpHW3ETAoRyTClJKeT6238z8XVMeMDR1/0bS2nFMKTuo862OBk
RDW1412nGfQLRYvgbvS58upfTCk00lQsckjJA2/IAXuqvWhVuuqVmaw2QI0y5qZEiZMg+LZF68S2
nSeAfniKGsrWrkloVSmfy/OFn8Q8ASies4tyCwV3sSQjbuTN2sJ4pnZkeeQBn6PEAwOgJ+qMGL3X
KWP/0xnA2aJHPCkmxdxnrpJgmfP57IEvUHeBxOIVXAxn8bomIucJYUfYSs05sLVMo2DmbHpg/C5N
z9QgQB3sbAF8Zh4Iha/XiGThlnBX18HsobZDvXsOtyiu2fvSO7DW2LxgxjaUi1LHQPnHj0Ui45t9
BX03KMkorfmPtmDEVzlGzS1M1McnQs8qNN1ExI2k836+KvZPnmbbVWlzKS/8pbspilqTocc9jfix
VspbZNfzCpwfW9YmJyKnfbuH9lfGPuZHZLRZ4SnmB9/6ShZK7FG662QMu2E4RXC4SGhDe9VInAIp
BqffHF8mllAZXdYytTEMv7VKqol2MPNqVC4w+/D842vr3zmnSAXn+tnHPlBIN5BVV3McuUtz6++U
e328jtyF8MMaMT33hMEY8wpQKCXhSGV1BlfRvhms/R+MyY8rA5GoUZTmZ8edoRAJApCtp+S5+y3E
pLjx3NpNsh2z1A5Li2bDlI0cauoVO5Q/ooUaexhxX8HCAElfh6XHZPEgJzlIFeafZwaikMid0LWr
tg5aQ9/TYuDnO/+WZgOnGenzfDIdbH9EW+LsePgZY1luNlk2TdbUzE1UeudJ1Rc3ux7WSJ94mfhJ
4juUCedicmRLYQR+XcUEx6PLmaw/TbYIQc6shE+83XLXE9rtlgcHz3l+ji2zsPnJpyZIyvRn/IF6
DKQM2iGEKhKueUdElpicVbsmISzoeANNrJfKBnjNPAnLsY6aMChTS9MPiNGMVC5RKgHosJDPw1Ix
PZPA5aPjVQ2ul+LzBDOnhbNXsdUxm80WHXmb1GTF98XA2l17vO9g/W+2t4FS/Qr0cEB7CGT87NP5
uYVuxMYtl06zY/Kpwfd5FVzorqK80orhP+2CDHRNQGc7viuYITXT5QpNWqKtH8a2VE1kFGQnKb5y
NqrNEvWhYy3I5k1rsEIl1BH2ayWPuDoKOSDIGrSrRedq61nmBaDzDoMI+XsWoKDCoYvmZubnQ5os
rDfFKk7L84tCnQwCfpG5C6MMSJFdzWiRw/3GF5BCX4CNH0d9SB4rBNFOtZwei2dlBLBuePbwK/GU
oLIc6AFoFs8SHC48+gfI9hbqPaApl0iyKWH5qEx7qeGSDnvDFFWvlppKqdocwO62PJMOIDv24eRL
w/9kMsLbmMmLc42hIfKyaIGzPUzNRR/SNDbcVhcPkFxGW1OW52O6OO4Z5SNBsgdGwF824KchBm+8
pj+6UtJC3Ov/bif/40yjQJhF8+LfUcronH7iFWhQX1+QW7xuulmGnBjo3aFrUf+NpIyRDk1dIOAv
xin3rI4rXBraO4Qhx8gq2grRtudCwWi0iTNwywYEyqRxeHq9HVFHzv95AA9Y60r7WCB25rAsv415
MoHZNZ6kgr8usqEUyjBThBq8mA9Vxbe5Mz+/NuMd55hRjn0Row0HuMESzHPzhJwxhG7ZNMnYTzFU
Z23pP90B61fntA/RWYhTrDLPCqVIxiq4KhURZdWAWedPdSHv218r9JcgcssHgoa2qUr8d5o7Ag4R
7bcICehsKKOmIQPMzw8b1OiMaMhhgyuRoYr3SwzEXVubyEOOO+UUIKaDAocdxv+s0y39LP8Cowzq
tc4ojELwvakpvi1Vrep3mA/RGrV5qiH5Aug0zOxyb8hGVsXGqPsz6eCCQ0AeVLyKv2zlEYox0SO/
SCEmOuOY6vfI+QDVNB1I1q4CrXQm44aHmWenILxhY9FAIeldD4hL9+Pe/E1DHZgbBI/iEx0ExXov
/CwpV3779i95IYQhiAOiRNUO3MQj5vt9BykfQf0KQN+vmxX9nTWqtEzEYsw9CfZtmpyP1JmtlAxo
t9/C3AtCCHccwuH0m4cYFS5xB+rsQgZNkl50VkBJZ2gDLqZ64pbJdbMjXDgC0EFjFpxu1+EyeETu
hcBXiVwtYciQ3/LJg5effm55nVbOjui2zjb4yzX9Z2QcJgBnVhAn99SDmhHyBfjYIXKPlG222iR1
5ubehuPKr7guf+XN4nkMMGLhXFY19mHmuudJkxYCUGzDC0RtkMQXxkKEJqAjqNogKSrvigrc0ujh
DHsYUlIMQRT6w0JSo8+fURBDThgsLZYARj51gA3n3mGW0Qkghd6clx6lEUCFrMt6tctguDQUsOXH
S9mFFo3V/wKUxg13RfPitIWFjey2zKGZtGfy1SyTIoU2Duk/FywNC1yZDa0ZqW/d6WfADNK7/APi
tLbEvA+G9rmTYeNK/KkipZ6CPdDHr+Vo5lmfL5szdcQ+y21YUxAsirQ5SBEZGzsn8Brtj+nP57AD
3A1tbAXchoLW2N80feaf+cbyW5a/eLBoA3xueQJA3nVX/3Cy8wg/ghqrh4bvjVrE0Yb3EotIRWqG
w3BSmTPCFPwGCdyA+9JvGwOcigWwj6V3a1zKvvTlom6JUPoU1K8srArmsKYuKX6e5vaGJUfSUVQ2
cQl3dPv7PLdoPG7tkb9jUom8K++eOBPDf3gOpLNksZiQvOneua+dU92SlaVGqaDmU2ID4HsWDaj4
IQstO1M/myaFAu1wmocYCK+809RA45JjiwxBXw0qgB6phjr9/CN4WzQ62BTc/DwAo90s7WhBf8ji
jvY/5gJ0OoqnIK7u3ZO1wLfRZOCv5phkMNgoUwVwApwziWlacYpZDqPlT1jNlXH4TKEGRrsmxWf9
gmWnNOUQMsrjs3es7n4San9+ZryHrz4owUdPE9XRci9yPaIbg2EcP22ApY9vaD+vufnXPcOZQsuq
1iYjs3vyvfF0zpUVxD/muU79xFTVWeuWWEzUwvn4jDPiC3k5aOkCGwYsiomXTrilJa4zrEMxZZZK
HIhatrY9QtsSnY1FpnlUbO1Zbyv7+0e1ATlPHwbljga+s1KXRGTv9JsVX58xLaUsoVe8eT/hw45N
5lniFjtVHuEWFFeFS7AhefXEwtI8hTWRD4yQEBZdOqXJzdR2CZko6yFVUL3+dZNCAEw9Wzy71CQ3
nIJapn814gQXjTN13mLr5GcwuvujWzakSM2iYrwlnQuQfgNS+5lWAOmFXuIqoH2JQ5eenwoyQTdK
T6DdE9iIYlHoFokaQdP2jalcB8hosSUNZ/YP+31e6m0rvZHO6ndZpsZEyS5jrdcrEmQoVzpyrIBc
X5f/kx9wEutisoD8pvA9vTZ83bBqbDpBmDKddkOdZ+HSYCjD0FHurAB+BfwAxSIMkHJYbE08TjKa
N+56Tz4SmayU1i+9tAte1HmgKjmR2w4Dma9LTanTgnwveTFHeaezsjtyUizkp5kwHWyVwtk0oU5B
0IifW0SXV8VoISMUVRS39J0J5z6THpzcdQe/DEmh+RVZbu9euEY/J3V/NPe37V2XBln3IZIcH9th
0+ohZ5dgUCfeGK+kUjwgizokGzRyPMIe/DvArC1xJK/KnVy4FTRsF1rz1egwNN3/vKpdAT2N72eh
7xA0VpQThGNOzn/DWdjr3UznxYjRU2+DtSpS1sByO59tqsKifhpJQgllAEK3mF/ohydRYM0iv6Hr
9CjjGftJOUoNz+eg/Fw0icgRK7ql7Wtf8Ieu8MylHqBs623dlbUOWH6mNjR5CdcmVKUPN4uUEYEh
ddNijevIlz4pz+PEX6OTuH0yhTB2B77sJz6HkvM/bRNoKmg3UryGebEzyDOwm+tpiTkMhwSkgGhd
l7DD38kH5L1mBGoFQhslKmknVOZSsZNQPqMjhuzBrVTNhHjXjozs62uJ4vWWFFlT0wJrE4gBkqu9
5AsVa76lTeUbEfzNo7110uopj2+X3XXXR/VZBg8TekACu6DuWPoDrZueL9Csf4wrZ2G47ayK2Lw7
P82VuaBk/cEK4mWqG4ejhLvWK+yC0kd0dQu34zRF1V7Ac/qPFq8RVgZFkg3v3j+c/kr3B6TSMxBa
KF5CvBefUu3Eo7iVTHJDGIFAoM22uluFD9PUMOV6Nrm2FZ4gY/3HNDAuJ1xYktUBLhX1g9aaLZ4V
N44Vs8I7fVvsVHdaGtEou248G160nmXqvTa7HQAVQ2rxpMI1kkeVzo/uCBDS6GyzFnzrsEp4Zlw9
Z2DS/OXqicqZwVv9Y5G3dJItx+cqVbref8UBIixgEdFRBirIWcw/c7ZnTAMsC2HIR/bTV/S7Mz+j
JWGZVU6s2bqpzvlq9MaCz3gB8VimDmLIUrAGFxGcLdT3xCKIppsjgsTYjjbI6cO+ffw4QV+5rHS4
eYQbRfzsCvkhv0fLLzletsGxDdpF/RTKhVrpxqhJiPTvSmVk/lPvwHRPzoXdMqSV2mczMXRVCcHP
GuurKxg0jXgKzi3D/8H+i9fhjhlOjN1GbQLIAkVXfnvWfAWZBrJp3wXl0llSZv7/fcDlPoKkKiyS
6e4FbS+q9p0lnh7WiI5OlpUaX9v4Fp5ZjoqQkk7MjS7fdWXwbtIAk+jOZSXILBMjb50Sh2MZQt6t
OPuySXy9AdMKp7i6KHPlgs5IxY1QvAkk6suznrG278aVQtTOUunATAd12OfnN0nm2R0YNso+vpPi
rIv+vhOKp1++dJCaanl7it/Fkgta/TJNRhf1lCQbaM7zMz34UAFSsfX0YlV/IhtzCCfG0Rdm2DB8
Q1A+U2vQEill4SUmk+PU1SNrZu/uVfoNEicr9pBfVRHNYVzCt0iLkuUawb2nH8BrojHrhUW5YKuK
LtBv4bXMGWaq/BxlqaZwddjEyiaJBapZIq2WBjHtdPe+J8hbXVjbty04lI2RQFBdyPpFByGOFtNK
ULAzK09cMT678mYdceNXk3Qze/bYF2E52b+wi0s+VuZ/68jvqSSBdgNcL4gYVVDoy4svUT9wpG44
jWBrQVcxhnNmtMpdYQ9XUBfdKOxtlcVNHmKdZab/aYUl8GlWQKzDu8m7hW7aqy8BGX5VHt6HaTd9
oBduhacoLsY19s3uJdNoCYgGkOHX68ziLP7FzPAhDcL0m2cpgYmwF0cNpI5yWC0UBdVGZYGb5TNf
+uv3Mt9oS8+YJ+wTw6kvt63Oxe5qsbMd/4+Azy4A9vepXiusYtgQipCOLvR/dL9nGwetgDo2CFaM
XQGBnZzrF4yGMPYPNj+7pZRXlNqSxVgrtS7aZf4bqTXBImHno3Owt5CXaOrlvhNHvGqVyEAdlVod
Iwp/ucxaLxmrA7UnKmUe1FxJaAhjbCQOOkRe4KCa+sjI6LmjDLOYLT+zwSnEBW1aOvP4R8EubMNf
UP1rS4a3I51qG68kNgaVxmZdxLlQd6L8LT0f+6IAqpsPn8UN2GIXGxAZDCa1rGI7llV6gmz50Ue7
QFV5GMct028uIfD669RibP2VYvlNYGYErcAFltXYeUoeZRcLLKivPYBBAcnIGcduwvyRV15Ru98z
HdZtpqK/DyB8sVtHMWKAwZK/0V3few3rN5ypzMBMIWBKR5FHgPwHUJCxTd0VlD6yaYG+KLlfEztb
RBmCtB+yJHuBf2I9YgOG4mU3Latl01HX3h9n0uGRWcd6Jp7396lqZhJgSHEUSdR2+wF+DHr03Sad
YIWrJFX3khHCq5G4sthcUxIXFnKFdxpfxLX6EKQ+2grUNo8m/dhooK8gU7MMExkQOWK/2szh/Es7
gsgpIuqsKU6MpuV5+Juu/dK4xbIac8c6OSXyEQgtNHEi95es2yePBFHtHHZo3Y3Qe/VIc1nuzPXL
UgavdYObv0sjZ4VUKWECyi5pHAZ1OoBw3T8e6JbshNZN4HpmFzWzEEsk0prYi4Agenct/KQpUsSg
umYOKn2PmioFc2dOUguPI6geWXSKe7w5M3GOCdVBJ60kmSeKfwop/tUP063yc8yrGyp+OSifJ0O5
WnKVXsXdeo8oQBR6jU5XttFsBQwLT+jHLPWRf5Wt3SUZctTT0kAsG5I90L26pq83lsdFH2+cFpGJ
oZ06Utl0JEqnvFHLHzr19oVtzcOMl0zDzzuH3pvf5U8XZfCdFzZm68CfpRXTXJxLkwOJ2UZdJKjs
MxUr3a+6IuonrP9QYfK2ZBOdKYAtwUcxXyiarkcFhwPerUhjk4aqyQhv12ga9aDoExPX9ZYZD6Vs
i2CYgGk8JbTj0aLD08CAca8bY0pUfKfyob4FfB37PumL7/SzTaryLX0xw/4m7KlxmyaD5qY5R/DR
DwIBkgN4D4Gb6TLKH8AoxfAeY9/C4mWURH9RGrcbS6SY4aOgzCIOattPp6f3GI2n/z6jSjwtKS3q
jgR64ZB7Edx2dmXfT9zENLvfegjXPaX2l4xBrG+UEqLotUv+AimI4Z7kIFU+ENMiUfzOyD+grv/a
m/2KAB3EewWe1f5YfBBC1E01zo44Xt62bETwpwCsFbPWchgtV8I1Ij0fJCJ+aF6XMbL4H42rku/v
Iaiusq6rW9QR7GGaN1t9Gj/1B1X/M1O5VNeJ9pcbl0CGfuxdFJTqr6NuhiZzDEdWLQLnR2lXmhi1
oTDJVK8x4ngf9RW0RR/Udsc7GYD8YsH4sa9v6n9B6FNwn/t+f2Jw1CYcb1fqMbsfDyCEnfT+WlyV
i2gr74w3THyXyJrkFkqcFKEKjhf7xQAr2ZgHHW7EcG+mbjyzVeI+Qu38BA0ekLWXDvk7UoO9sybN
OT9syDyyIjUcX3dIozMZ5GgwJsaDjdzcwS902u9VPR8OdZo8gB61/lBGrqgbxv1n3LcDXr5WiGJ6
sv+8pWtM/OIoKyWgKmvJArjUdSAdKKnkHOhfAsgVqPHLY34Ckar4tptYLuwWmfiY8LaMAUes5nF8
v2FVYb9rAJoZeijTsZFeRq4BjaGCQon7GV5m4Bonx4OdlMOFt7Hwx/qbT08UwgqbMXMfTkx3AZB/
XjdfvYX9aGJhOK9obY4rpbCaMa2rm+xXyJEO+A4jlz22m3IRettFNKOnDOrZrYju1ZMFDu+zaJo1
pgg6osTfjDXloOMx+uXiPI/IYIYhNO7vhm/oVzmzdK8wZMv2Wv9xweL/ppysdqImkUAU+FwIpI/d
3zdu6XAnUVlXMEg3F3aUO0WL+OfdNfzztl9I3LvX3GVcJZpvIlddtkwaTt6PoIAyqHEcsILI6YcX
AgZD0IxQRJ06QbffxA4chmu18FnNU2IvLJQw1XmY89Agfoa6KFaGBhueAC2xuKJhhrILDLLlKiVe
Pzgrvm224uO8Tr4YI3MCEbTS4tRSq3ZFYmehpsspwAYNBiFQruuWP8X7LwBTTdrfwjGOZ0HYbM7I
puUaDLfE5CpZoYVlOiADfqcMjPLPEmNziGzG+JZ2Rp/h/y4NmSMZ89PGURc9SfVYueoP+0u1EDsl
OeCSctMwlcvCjLjZ4zoIWlHP+su/cVy6LGHYDexl6bibGcqUCgvU9ng+huR8Ek0GMibFbDaP/h8j
6AEL/p1MhvpDzraoL65frpZkalb7VjerM5kXs3ziMTgC0JRR2Hw8X4FcsU6tkKZKv09zkMhv837r
zpGd4uuAkK6rRw7CP3+zluTAD/77UtM7UrhejX1ntAV79esdHVL8xoK2X7JMSBHATMMquHW2UIv1
5yL1EODGlAIh6U2nREPWxbPOemSpNp5yGsbZk486hmy0WUgLrHGBYUszfvNTEWpNh4NOWoQrVqIo
ihYeF5LXU9CNtUBwcz40lK3uK6q7u/vjs6dJfGDY9Zeym9+Za9zvZ0aCFjGnYoxMr2ZGAsLBJx3D
kGKvtTA783DrJtPSjLfhvjPUJIp55ctTnEs3yCcylUeZYE3gMP40jEY1yWe5CCBs00TsVzcP8Fw5
XM8qgUEVo4Sr1qKH8SAMuckW429p0vPGPoWgC+dIy9JlNR+Yri2qzHEp1kYhaPV8vIErCqlHGNvR
MGlOXWz5v95SFDjibdOGRB4RhS4fcFLhRd9oGQttfrjBe/bu30FCv4hucR4bXTb9AgGAx1S07mWp
eVRGg+ifimxjL6SpfvpS318wndHb2Wc1x7I4RRua1VBy2JpzM1DZwUt+krLi7lttr05mq60RaM0G
5tYAbYiKrMMokcMnHw3F0acEEuDXnxM9kh2ligeIBkf9Fl9O8imK/9yXWiVeYg9sg8Lbz6bT/K5J
UvBzumMxDfucKdVBDmDh+IQEfGE2dBADGlkzt/XsR9eQxiWcdVZ+otN+42MlR8gVcWZZ+GBKmmT/
Y+xaEUYmp4auVZZv2/UL3VRl2lslDm/17H3PJ2Im3lXeZf9gRf/GQ9/Dr/FAUTZrUIwKrD28HVcG
N6oxXnuQNESC3tXRQMxUZhKnv1nieHZOIvhGh+KcKM7JdoFOSAHSMK0RJ1mK0Fux1usNADt7gaXm
AJwbAgRERe5pXX38//K+nlND1U4mZTWsirJuWbsEDZ8pe4p8x9iLSfH0CQbLlwl+tm0dfFRSsQdT
gyTKpDpX2MLBqit488A32yqXWgThzqFXT9gHAxN9nkH0L5dXzL3LHwrZ2BewPwStvuN7itzIurrN
sP577EArjBX/dyYj++xKA6B8eVtWI9XTkxF03tV3GEXRPmXc9n58mkMuSv9gD1Jgz4zA32FyNuZd
DRMdOFuS/B8niSVdCcSdUQSAoUnA7NMIla5U0P4567/qy3oLuE3sJkd6cnzoNRN4TRmiR9cMvEmI
BQhBhftVYtAfFVJUmdD8Jm8P2W3gH+o8657DZXSIJWzkSXxmSA6UmmHogATNq6s7a7emsGDA9Epp
1+eF6hKVPxbs32xnovdYbdz5cpkWV1ehM1p6mcgIhuYpuRucQWjkw64jKhonOJIGnrTGclwwVG6K
jNKY052zrPizPKXDnNPEs5SDW/GciTFSQUoR4ApYiaMKWkWdldd9ZTFRrN6hIWhlG/auVZYFv9zn
8djUsXzR+aH6KFwCcqWfZIfukKs5opfXulG8PscqY/qHNWSEgtUgwQn0XgvAt9YvP9Aqmsm1nh3A
Op8c4w8cHpg4aoz1w3SNfgdNzCvSJveTn7cKjyvgLullS7BZWBpTNNkUk1RsbIw/Kojrgo9Ei9z8
BYic/7YmVBwy0fd9N2yJhg4qn93gmcVtzRnrXj1nH6ka6QxarFLGWXYgs0W9YL+vJSfbbJ07Z72S
vFrTiQON1S1TCXhGaNH27HU5pSPwKiqlH0o7IbJa12VYnvWH+Uac3+CYMR+utDmosdXmJnsqGe76
49fj9kt7A0T+IHhgoW4vQpCWDhx5gKp8Mu/+JyQtgE8BC5N6ricpGGlVpdKeab+1GqOrI3wO8eeE
QSuOMBwa4fEdPtKqTzfIZE9ooHGC4WXdHtYyptIh6o9saC+c/BrWUo9wzHfUcVTwn9ml0P7UUGvY
p/6pptkSCI1GX5IYXfPfzJAACd5z/pbqG2KzRwG9JuGhHvkvs5zp8CLX8OUZ3iZ9RAUEjHaohhtm
BzVE4ysLki5SWTJB/Xh4eRi/rJIX0tlJa2E7G71+bOvrBGM3qiq66AnjBqVnNU597KvtWyfN7wx3
7k1nL9jjxRA5RJ0AdlkDyawKZARR5i5NmgOAVXVm5g6Qy0e9zOBcFctYS+sA5VDq86+NPlp4/RjU
UAZ3cGWcdszAAk8BbbplArjadqepNgnjSMYAImEoIRCiX/+TvAmPSGa2B7UfFzp7Qd71LHG+3fyy
Gb89+vFmp4XOkqnd9CbinN8sZWjkvR/h9ocOuiWQ7JdyRaqFy0ZCD8wPmA+BN/abT1bduOdefTVy
11EIc5is7S0uAXR45g85hc9LugjC3ufkZfVB+CylIkR8VwrgPbQ4LM6S8BMFNwkpuzxwdKuOOTGm
B4a3eHb3RuGzw+u+HnEAuH0zeayYbhvhLeIExWgMLhliwp1C4FE2jg99kE7KIN0nbbLfWJtIMDT/
cFh/W/4x+cUdy4jqWP6pbbxzEtrNGeL3mClKVcnnoQrVHLi3CyJgq8OxUBf201W/hH4YSNipsIb9
jS7MaJ4mHrXMiHAMLV4ymaCE0FKXSpoB0rDeHDKpj5Ok85ucrj3zdD0ci21V4bOJPjnOm5ktxYOM
foJ3veiSrXAJdjm7ZksD97BJkoPvAdkbOt5xF1jrkXANgyNCdw81YiZ2bo2PtBnrZteBwYSXWrN4
Jmm46o3EOf4xJwsfRuVMPgLJ0YF8Ay1PgJ8NbXRq/5JQnMX5sRnGcoXSdc7zUHb3kPOrJZtkipqW
aA/u+Z0cekHBU3E25IV/GGG1ArYdlymUkEx5qMzGeEBgNvMftsZt20NKZobjRtZaRkYtWFmlDNFG
ygYfDvuOdSqEV2//7R+NH8yZKY7ED6WSTKjbh/7+7WnSXREV9MBsRF9K9+/+VnVnttUyJH3hrNya
zr05KNhtA+wH2a8t0d+w2Az6R+pm1pVoUK70JYZdyKXwkzZ2JqXUTk0L8gVzmj7pU/11niIrTDrQ
veDpp5VAP0hQjivmeUUzoCbBeFhUBY885Xa2TfBskqAi+Uvcqw1o0BmBFuR1uKy73R6vfyDXN5FC
azYl2UksD3lA7Wv2WkqWpIQIuXVRXVpXEMSm4xPRWgdSF0A9J0RigvrXNNzalNfN3/yQuvWPnQs8
oWvJMF4sw+oQM6sHn96ZPdVdCxRUIStDJmEb9TgnRtPIKSUMq+4SwBGx9xpabbQg+ZPoBfTXR7tG
+pspNYv8XZP72cgGwHyL2Rfsm2LA8npXDtUkMBWfYEFtlBDufh4EvZkc3DeK4rije5lhH/PXLSdF
8nT8sQdlhr0ujM2zTy7nze8lRHxp+Wesrygmv9zfULQA1L8a3GUabTo8tqm3pdcd6kqbQtnEJgpk
jKG198NtoeggZgYd2YYTLMz1hQijXPB9LI5bqisfsIrF8Y6blakUqosZC2lE/7GmZbAi2xeyEF0w
OXZfHL+H9B29YkoXK5boglR75KwB1bOcQ4kZia74rN0O1dU7nsfhJlLFwWjHzBWp79yQhrbYwAtT
2yx6x79HIuZkQTVCqOU5OUX5LTdOuoUVcV8WTfCdSYazYlMO5YqQR/XLLf549Iw6W/ijajvgUgIp
PTASelwp/WKk7nEdt63h3+dxv0iY4F/ivKY1HS+3Vk89f3mw0K9s8Aq02IfnMoqK64Rf65Rq2R2a
T8tseMQbrlrwhox/PYCfCRnXlmiDrhaXYU+w2wPsFKwNkpHYXt/tkJPYtXEP20JPyNtJBFMTSmwZ
77cqCKORNDNsyvhC3k02rfyIB676P8Kj4TOwUn7GGxpNzH2yYdYYDh0aS4sg1fla9WRXvsQbDpev
SmaqzuSPLF8xEbhLMY+xeQHY8KlmaEp3ph0Ud65xzEYnCpN5Mmn9BEw2NbequRCD6hAPYE9xhwsS
H1AKu6kvkzQZReOGKZJPpPT/xK+fL2rE6K42HzpkGJyC5ZfJZRCq8b1doC+IEcq41gN9kFP+2+r0
e914hLcApBRHiND88hpgCvweL+sy6PZLetH+ID900o4bL+XAKSHyTpboC8A8LFwO3NGlt0u7veQZ
MEDcyBXTyZMWnya2Jf4qac03sflNBFHOQGbCBUutp9Y06+YfqT6IeLn4YGrHuRHrDchnfS1zQ6YW
Zj5+wHzq7MOdpr4FnXxMN6Bzuq0kJR8B8j6vJ/3hb57FWpuKRKwhjxcNblCR3OALneb8+cddpoc9
O6J5sk1v985gAlGzavWC0XqmpJjFIeGiH+j8al3uhIzshzrC4ExwYhcX8qYvNLK2st5B3sZ047lx
P5JhDKXZwJ/Dl1r4HtuNJyn+l3XmDCesXOc3DIaF0yC35/UYep0EhGD3w+T8Bt+ksLb5qVr1j3yv
vytXsH/dtUOjT+AUtqj7kmVODH88hJ3LTAFI24ee01bvsSF1awC9u9P93OIO6s4CRBeDhiVwg4LR
iWq/Et6cpcW2nue4WTLcidJzmO6LUyVlgP4IR9H4pnSud/VP3tFO9g8G33GJ1qRg8bV3/6DfzJzb
lun2Yptxwll/jroRwps/wZLc4vEOaUXUcxd8th8rRX3Xqrvs6CKwo6rnhT+09laz8q0oUgphO93s
GTZLxTJNw53tuh+98uSUJ3CNqjvk19X+JJNTBAFU+hwOC2VLsehG1/R61uFDecf5X4pHdFK+qHw2
ArXw0YjVkBhUwmMhd1vAXWBIQhi7YpT2NAD0/cKZgiLjOcJt9QlvMUUvJnXHy3o0lwVrCf176+Ta
gLngtn+uAU68lNIWIXRpQHVHhO1LrUtpgd8eN5yKUaWUw+Yvfme4gKoEC2uBuGJqvgRGILq2TOVk
ednPMONw7cn5GXMftMSwhcf/IIye8E62FnOc2EbPDIjsJ6wl5Zk9A5H0TKTfmeWn04CD8f/jA5qT
K/CDjjqx06WKF0i8Ui83Hak5g2pQZyj/toODi+JyiZlcKHf7uz7fKXjY+6eXP0yJNfmMALB4XAHO
ZBF0jI2DbkWAAScyTmC2p97Bumvb7rIDw49AxliVr5N5TP4KLV9rkVjmJ6TdwQgBnaWmDvZBjqRd
H02MxJo6NTaokUSc1kjQIuwv0gnwcxrCPx5WhhV/jU8992pDuE0FTcH0sLiaUrmvhgiJrJXyphbw
OTdXwJxzuLOjwIg0tD6V00SOJvQR/8/kFztJB7lRfxIldALFJlBem2RndgpQTFwhvJAM3vM2RmdG
I3ZGk4E83Py+YK7cFRwruyLmNSLcmiGLgJxOYe0k1NtqmFGK5Su37gPUQB+E8XZfGyLhOz9Hm9VE
GW5YHj4L24NZnQEu0db+5rC9dTSgnVxQazFsLb7IRHbFaJJol2Qg87LbEVGjIoL+tW6Ww4Dzh9Xm
C2v48U8N9MLcl9Csn0O9b9UdGDZ8pavOTvcG0tm2xEeClBwML2u/dSn0Nj+/z5jbUGPC8A5+HyIg
ZxYwKT94Qgz6PV0LZzAUk9udrXEaeUr/bEEJ3T6l/7DCy/nJyfL/cnJ8VNDsmEz34+Av9qg8WroT
/HOnRfOWKyQ9QWapRBXnpNTE31Bt6ixvJo8L2+9QpQ5Cg1Ag5G42JZCHhq7vpO1isICnmcr7rZAD
OUOrciGaQHwlCCALc24yv45oPwscJufxyLfKZ0RxtIRKCoT3AKXeEa/cuEnzegL0XF3gOPjoek1o
S7tdLrFqr3NGTJ4ytdcGWbeIi2UU2+G6FjSCyOnyAcdXjPpLaE2ImwK2pU9rjY492OQI2k6Qn3kI
C94lFmq2Wt3/0EFJA6bZvLB2uPGXpeAQ/13XEJJKYmHVE7aioSGGGztdgZzN2Ydw57NrQnYxx8Hh
E6JyWVTCPRM1OR1WUmy1tTli7uIkO8C5BDXVfHmy63U+/n8QSkmxlgOCV8NO57ryWOz46y9wAuVN
6yr2yLA0W6bBGyFDy7SXYslMFKGCXkEIlupXcDyPwW4QsPU/JceT0nADcG+R2Zp02I2FlJOfuAXm
3PSiZagXylZ6mBFCwWJajAzT9dTb6k7EkSxLkgiQMRo5/4Fj80R2QZCP9Sf70wZ7CGe7OxjE9j5f
PFkNXubg+EN8Qo02ekNraH6CvAdy30jnyy+Uprwk1YhVYFYRLceqOrI7+xshg5s6eFM4/z167v+G
5eY4uehc60KUJ/Uy7qWlrrfWf/TjM6nGHUjuP8m8F52MNnVirl4AZ4q3YZdnGGyU/tPIMlPrLuU0
8IHHQwj7F89SmrOPeP1BMdRbXoJk5MU5ErvSPeJ3svCCf9UtIdqJGDhm25h36JJl9wQh9NOWbiqe
AD+kvAIGYEPt+iCdNmQyNfCvGOFqT8UWMAxFf6Wz+oGQtNiYS2tb4UZzpV1PtIgKfwxuO0VixIuV
erGhntJ+Irrz0E7aZmA14nlIQ6A5dGhNc5/qRmJkn/AqO1MNzwRQHfC3h25EtDyhOrCssr96TTJe
UIJTWITGBrGcmWBE9ixslephUz+4NYwJtzPsUwkMzAdzTN6qwfnwRhBvmdKu+umgFcDWycnbSCxh
7VkyU5qyXlVfg8k/gqtxfnmnQp0GZgB3bukCzWzJruRe3GZNcP0ENZwb3AlNkSGqy3b9QFZqnzGB
vKeEA50xOZoFzTKIy66qdYyBlT8c0OMbhSAZDYomtUPjv9RZCwXfjircByebws7rhxP+F3ZbsIjd
j8GU+MEdzF9FLvbCZ2DDcQnUxl/681QT9KC3+0zeBp+MjD5fSAQHQtUxah8pj/AQ/CYJOfpdnbhN
UUpXKXIEyV0QKSC2W5Ot5WO/8MQsaU33g0k/mqrxzdKUvd9xQ4HzY9m0shyFAueny2XQS8SVvus8
DCCUdpgNubzJSw4nYlG/UPYDM4T9tfyHT7R18hbEKbdSptjVYlKmLvP768kNv5y9G0TEgLsJFIJp
y0Bbrl3jzWtyYutsnoPWMS3uigwJab4mqbwfLtXvhBLcWYr7qVD0YLPUSwUUS5aG3tz2SaPnujO7
24xCTeVBkIkTjG8DI4lUPkhj3IL+JGi3xF2sWMjBBdJIEENHZsth1382nRDAIkr3fBsV4cBIXMJi
uTMszghHmR1BQ6dwdXv+9xnwyjzMuGxkpmDiOWDt4rAI2XyBOiQiIvpcjbiJAcXsmc06mdPXiNxm
kaV/OYlCnHYWYe5dpJuIdKZS0ufwxhnGfrc2FozbhnlPMY8YMEFLkjIgA9lTCFy+Z+NyDD6pndqx
t8F4qPr3WJAyy293hkJiWzW1lF7ckToayQsJMSWis9Ccd9C8K2LiXNulQs7z8vhnyOwKGvrsgLpl
6caOpxSwVJha3uzQm0yz0D8mn5ndaqmye4dlJSWLSClgoIeikAb/h1xYP9EFmQjH9FandUcwTzMj
wD4yJBTJ5bh3DmyWcxCISaKh/XzY6fJhzHyTo9ARq5o0siS9eeLGqIxpzb/tYhvZyb2bPewu1vbc
JoE9JDAp7KGlcjarMA7RCUcSQpNlAc0x5qYxz8J+vaRXR6RjwqPCh+sD1nwTna6BspZoQBWsb2ck
E1kB40sZ4o+0uEF+EYZnbbva16eEy32cY7PJ5YkRBjTcOXfMnrUwuljVRhtihJ41FFNJFAH+rGV/
ehnXiLrS37wo44zsxN12w8gaxRRXZkJRhHc+bYBWOrhIruIm3+R/K38YtUGxK+ofZzB2PoGjcXSK
M/ZeBvw65P6wG4JWm2sipAFo7mmUOevDZsxVTZ74jAUoS0y0dw8e0tpHOnEu475R8aPhrNkiKSry
+EZJjeVVlkbpgSntnvtlOfBSgOI9ty10ILCdOExDDkzu9Rcixim8LmtKw9Wv7blyaAGyx91oy0xC
ZC52gwp44o/Yi5wPe0n3ngu8ncB90u0ioe2qT5YoOL7/IWTMBfo0ukNVL5JJWQqRX5V4pJ1hUyGw
JhioJ+ywx5MpuzZCCNEgzj/50FAwwDOseonzHp4GzDtG6WSFX8zJolg8cT1v7gAHaLub8Fq1iAqN
d381mykmss26XcWmoU9D+go6+ddFx8ukNK1R30AAuDnRB8rgxtMTgBzr4OmWqmhyn+WosQN3+ZGF
Z+SvENfh0fJ6DeqWvucEMT3Fp9G1OqCAUQV90RmSUDd/9ahFpbzk4H0KJbKddSpj2Qd5g1YaJlfd
z4z/EHzN+SYK8S4Y1cyDvx6HN8Vxl2ndWDHUhBOIaq5qSgF3yaUkIy+InJCg9bex3w5DFvRUnRPz
/xFJjhKsCqeoZXVV/s4diAOWqQ7sh99KqMXVI+iTFwZww72q/mbwFybI9MqV6hs56DIXLl+Gvv7e
ukUqZwgUSm3hHAWmAgOD51SkzYSEsVAdusodm9yVYG3CeJQWBSEby10pd5WhgSTlhEhnAV3e2XlH
igtdBFhAvI+EEykTbtwzcC6Rk8HClZhecf5Dw2QylCi5XeYiQ1I46NTN2PzoZZ0RZbpRVWa6PF19
WbtycKZpp2a9A1C0glANh259Rd9XOLoujW4axfwZdffeuzXfpDvbwJGVmZfYG6bITJHLoRjxsS1c
woNL0QxvJrEKSQzzUarqDXiukwzTe1NxkaIAJzIvaH/Vp17F4fdvngCkYMIpE/HrUFu9Wec5xCI5
1ceD6WK587wChvM1oJzpUxp50KQt5IcJUt6IZABuAIPewXOiwsR0tzJzP57Snr7WLgnPdsGaHBcs
lEak+nvQLKBZiJBuvsW/sVMOPmfx/AJJbeGeoMty2V1sDeluVoCdCz/WnfzDxTpYFw3YP953PZSi
YkS/DAFhQ1cW4rrkW4L2QwMMeDKJbEzz1bVe8FtGIMWq0jiNACurch1DhHuOCF37JZZmx1vPSvNv
N9bSKHx7X4Hd3OYF3wCaM8bjMVETZQwWMCCSOCwLik8Vjv9UBvjuc1E+9iuNMmLWGi7qaOGLH/so
TbucFanO5phuWhMjBcxUTVCna8bHKbLGc20jo55SyPCWa685Kn6U5ZDTjOua84+4maoUXHGDKLyy
lQUpArjmLJtnCj5nJkO+smqz1vyKsJOuULEDceQdWLtnGmy2+DGZRdoYxiOSzttl+4M68XFfn9aa
zXWJQQLZLhk69txCxTbTPOmmghpRQoeidHj2JHnf5DjtYBwdqbe2x/DIR7k9PRncQD7PKiAPjYoi
UFvrIFAzmdNQKvhqrTsWxuzMftUn2yias+xYr/ARu4c3qRe17j26fpXZ+L13fbRIP/qNdimkEyAD
wudNxx3LI/z8HouTC+mDk0TWiyawOSs/xcRmisUh65mNt3UsLkZz6IWdsouianZyLKUWeye/N/SY
WO6XDvb5k35ltP5E1w845bk0nnZCQfgRbiect1QGs/2UUWxDhbJJuoj9IZv1ulmKCLXIg8uDMOY0
JCQagGwxZKLNOXQxg0Wdmzh3tUNHp91xmRvme8f5qn7LA/EKXfL2uVLwSlCjaiOEJKTQtlWGgtG9
lSfyIlCK4roDuHIFfTjn4IBqu+3eWDJkIXe1NoiDeYM7RGASwRi5qcDXtwx2T7JpM8SXqrqrbRVC
++3KP+vlnUHs/l1ZlNM+vZMIYePcIyPL6KP7dcE+o55sUwrW2Ipy1TazvuR9vZEAPticy49waKhl
TqZHYfze0wYsY7aSe3g1e2fferxOeZ/qSQGVY+wh+OnxHPsfAeJh2D4zmJ8s6c4cTHIA3jWtUwfc
dfaM6RCHy8ngn5oYoXmJjT4lZgXAqnniCLzWbPsrfKkyRp7NXm8jXgooyYJI9aOljL5KqV9quCvG
lb/vZMsWa6oMGwDvq8jp7tigOiomhLZhpX198+ezrHHMhub/O/rlSvOsdvq1w7Yks/9tjt7P5Pl4
UbMxyjwIsn6dZDV9ZoxMhJCfn0jQRT7dfMTC76XsBXxG5RGli447TygTHlvx4xg0bEr/RwSxHI/P
d+FrOZLGxuHY5fC1P188v3DA7/AZ9shotDMGeMCMDzPtyPxQE5fHDYOtSbn+pW46WzhZq1yQHEK9
wdGkoMafLSjI4iuXSYgJ3Ykqyi9Ej/EaMcPZSP1YsRCHrLUzMsjNxZrar3sq+XbbdOTE6uQilMEQ
QKmqmA5pLJK9n88LP2YNCU/B0ZkrcCaFf3LOJ/uFjSZ5s7IonHyP/MObDoMLCNRruJvXklbnV1Dt
qouZF6qJA8OJpCyJInWFeEaj8PQ7b6yhJFEKLZdKiYjVvQBhYc8IJIjCm0fEvTfiN2FtmX+ny/OX
BIo/HG0AKgENOA5JaBd7357WMcIeyL+LtbssOKl1pO0eWSRLK2ldjlquveQq4P7j81bkIs5PjxJk
1YwBbxwyGA6sRb8MSYePKFhyAjMaSaGkbWSn10K2ehDoahu/6GKaN16wSdCMQUvP49+vQutCx4kp
UuqDkXEVvScEWL6MGZxR0W1qeVUESEiHo4uFhP+yO5ESyEQVGVvOJ8ulXOeekkANxqjMuwRCPIvT
+vcifcQt5JrAIlHbC6rDPZOrR2Tfi+BaQN1NEby5/VZFaebQekjdl7ZzKQ3Nsu8MKBojZqdMLJKs
YjWy6p5peX+tsqsZ5X2GvaaP5GkueTrT9fkq15kMZCsDJXiSz+trOuXR2m3VhISTaJSSMSeZBjke
VeDZYCT2qU85L0HSs5ymMvQpKhvHBjJuB0+frYZ/+eTr62rCmJO8uGcKeFCPRDVb90pjfE43pBN6
lIppXT40e5P0PmvRdIw/sy6zQp7G51OuPLZK5HbMyyJHl52LdIPauZUBWc3px1S2wWLb1omxLLBR
FnSUHyWs/bhNCtyKW5XVv2sc/Bo7G4JLOeIZ5/8zZ7W3S247AfWCvQHaBZVv96k2CdDWnrzb7cLE
DL/YXxqbeGQYnz4+JtvrL/DgMFSgogqzf5i4HipZJDOyclAxeGyFW2tTxXz2XsagKFlh4M5tRwa0
Lp0OfXn6q5ODjsc6srsOzNCX6cnbfpOYTcLoIO9qMhaHUyvsx8AH95BShriceIjvjy0OVJIu+xWT
bIns/v7DIqqLDxtCJFgcdFlasIf4DTpW5agbvpbBfX4lKGnk1VePq87rI6GbWUZXMaqUyzg0xL94
Ng01wZ+Be7mlvYjVycnbzHB8Z6xho4WTieoXPjIGeXsalKxE7Y88PcyGDCAi+/DSXUwSg7oCWinE
OSWUaJpCJvbCTqcRs+ylXbjmiZThqFqqJh3bSbaG9+1JEhiaaTG8+xhO5g9Sgf80G8gABIuDlBps
WllOnqZCfLU6U/FiFC0+klGpYiJGnohBQpNUPMGxp5eckEGJ5CMQWTeOrFxq8fi99WSCSIGsZGRl
naI+F8opUIzsrgprrxZWakXJ7CN78ENAhd9xGsQQK4+wrM3EVN/rOlWyOkbtslZTBZ7IDbZkp61v
zmU1XyH2D09IjnBNLdmNJm9J1tEI75Hk6GXegmlgfkbdQkGXzZH+mCVknqlmcYNLFOkSfqgGvzB9
DCJQf0yMuyu+K4NuDJFVdAWbcdTBjlFl5rkLU1CrG+Whaj98EjFksSwhfpk856coRpDnDDET2Hiv
D212ZT22zEQQKP1oXGbfE+aopGPF0EOmR+BgAl4T7VYtBlLj0CXyVv8h+I8cjvvmuaUbIT0y0REF
+GRA/7Fekpcg5V8wFyh3nxBms5EVbfG+HDPJwbyhdyhrBHhTk9OrFFVX65ySes675+zOxtcUtGTz
RxJTo3njO6y17+DEQ17u1hyQ9XQhIKmf7/oKTMQrFaaSjun6z2UjH4JBgNaB1ENViEBpf1iPzzLe
lTeQAxmzrzavksgZjztNR84f5tEAIASPf+L+YOZOs3ErwYNZ1hZ0wfkfmnL9Mausie+DMt3qhRlx
yOlGi4fS4EnwTj8790gkldcMG6PAbDdmQWPLgctPoPAOycJOFg5PcPJlBblPC2hsU4UXOaBb3X++
yBsasTGvVb5xGuBu43jLPfePcmIXdIC4JUP9T7tKvwO8cbTto/mLzhJtfyU4OD3eEovxC93XeF/d
QNExyNnWanexjLJ8Ku/DOSX8fpSUP/Dld8PwCxJjSVpfOLd6C4DlkPvCC4I9TcMldCdM6A1SQlgj
ky/YRgI1/rAFF5QpkIe7v+Sj16RWSXThua/O5id6aGTA5FCT3m6LzNTezebvWvZpnXpWNgbwDTFR
yS2PBFCANdgzc9XuSm5Tk1S26BSLp+yZqjQX/Wk+uCFSHKll2vD6gBruYj4Vm5yNngrjPp/nPitY
CCVmAuR056ooASCUqfbURvvOu+bd0kBB/U9+VQG80AaM3SqQ5GBxbMp4OlGEKG/CDEPyl4uKtfTP
6VfSZlvbMVe62bG4d3fgBDtfzhCEuR7t/GC8anrMMSahsaTzgd7rlwr2GCBRL7InWH+W0X+Auci4
phCc53fWJTLwqqrnvMNOWaB19xAlzf3M6s0IPLKoRROPK2UvcY0svcPCpAh/gAEgXp1j5KB6WOvj
NfUtEsBYj0hftUUOvWi8/aLqNA/mbaFCDjH2bbGFl/Lgy36XzB6aHY+RzzJTjbaz5NrAnBdDe08f
eTqWeT9aIpbdrIKDNTphbziJy1HxDbeIUQWnhNFZ0FUMVKtjMyHPScdp8uP5MUF2j2Tm3I4y4r7x
WZqejEHXaPywCSyN8+Zl2VO+SFcAIkcOZKWaQWsKbp5VCScXR0swOq+2Hk7iyJMNKYTCxDMfqYpE
7cWK6FEDmI7QcdJlBuqF8xfPlRxVIp0UNx0JIYULv66CRCWsLqLbqksE1MWuuEbCZhn9uMWoXtSY
9116vj8EbWBGmAdSWS52z55dtZ1kezw+0ooiro/V1ELdc1SWEAdiUgULBGhPq5yBYZO6aW/UBxuz
cxMWp8MmlvYFlHhbClg3G2vmRm2g0IyJvBM4+1u2p+gT5cLnj4hS2PzNu8seLFPM1q7Xo4aphO05
BZMFpraob95IthL2J9LhRZZI3y/66lyeJ124jWW4s6vYmKI4tAe8A2I/VjsvXx7zvxFIFOobMWVm
qTDAhspDXaFQ0U3+x++kwCb4IanMkzSEZE2JcbYA/rFIt7RaXh0snm7jDplcwLSseLXHu38akrDI
70Tx89+s1rujfcHeznk0EeYNCBrMUrpvu/6kgvUJIxjojtfAii+oI2ErHS92eMjhtUbkjxLmgQ3I
ZUVhqhH7lAWaiMcYe2UMiz9xC1RSxHsdwSzlFXKdljnY3GrrckzE3Tj+O2nwcDRheBkOF1oaYki+
M9e388KcUpO6zc/rklUvQbZGf5REsNcN/FxaKBkm8F1Z/AvkoDBBkmkyueJfZAodiADiBSO5pmiC
iPbhq8klolgBnLwPZH7aRzKPXpEUEy/wWDGWLWGRou056ExJM/4jWdKv9XF3cZD7QNxnj7+FZDUE
yRCRoUVKfIv77eNMF+Zy2gP7FheW2kxrxJF/Aou4J/ZHmhMyOcikdAPRlU4p6TsgfHOHeZsq+OaV
R0UY202n4iDpoaHwRLCE02cJc27Xg4lke0SpXt+z/jyFzLPXtEymfvWy/SVfaUw1RQGuGqkhUkcX
5dafSn/xMtFtm5Ma/2z0OazyOO0iyEc5R6Rs46vKU0z6vz3khiAmYLrMVO2iZO+Fo5RgnYHv+QNk
eJMB3wwFzEAB4btcJNd/6pChvBQ35d9Lbvzxk2y8aFhhvbprKI28ocDQ3kDKgGGGOruQ8SFPvc/B
VFkKmB3q3ShV1HbooFutiDHganaq2aGAh87ndc16imvIqOBJPi0LzukusafzGY52WoCdXGjFb8Bl
6xUJOGpSEPPZDWOGQIo6IsCkC8UfS+daWvCr0EyGDQKHINL8p1oi9nGNirMbuu+vO4aiOHqZ7Xqq
FtqVcjOLo6/SI1brE7oV6F835A/vDI3X4yqQ7QxpLdO57mtDy6eKCV50RDKLN2t8A2Hw+457rII+
TROrBfHcoWsfWqh6zZy7cNB8ngT0rnHaMp6wIbj+EQnmUdbuFD7irYIXtApm59WzVf6kVBPZbc5H
fgMp9KQhEkJ5xruZf/YbtiNJB90+inSTCXRs+plUl0UfyN6rGOLnLHudXhe4jzWzbpWymecf2Xzg
EwhWwnI8ThiKE4/ef1C7T0v4NALjaAKJ+FxYJ0Q+YGXXZQbXqdUg9F9cmpAe+SV3bSrs+JGdXxDt
wHgomIRzqneZo4csAHsEdG1SzOhWPH8uEeqKgUI1aLUgQIwLNjyGsnuMi83WKAk0Kh/5NMY3slVz
8TS2r7hXjUQqcBx5OkhLce1nKcrlIM/1RVOAgtC1Y7WMZpWiIs505Gh1LZ1fGR1ox9Nf/H2rhRku
2Q5iuaRpQWN6zIc8D1r0rknN8MMG2CDHZwsottJK6eYRvdst41OS9b4j7J4qADjISX8n+ezwtnrO
GI65XFn9BGnGJ6KRzg5ew6mDj77n5THhxIA4kXaM6n/ui71kReUkBpcDXVaaIxnANAPXUgVDYQvg
40i9fGdO4T3VWmw1Q2ERnbGb2uwDZABW/qBUppyNkMB6Pwovb+bSYJh06TygjyXA65+Az4RMnynl
lxaXmgrpgTZqgzfx863fYZ6m9LBp1bcQm0R14ohMj//P58MdZ2239VuXDiW3VrHFS64nyefkjj3s
X6Vnxun1ydrEQSbrFb0S2b411uSvG7o0DuwynAE2Oi+wiACyvNBUF9YFvka7cKewjzMJnYM+wzLI
qoBuUplkv8mGvYgEc8oYEIi0fDJViWZhwhG377oAbF4s+tlQ1/E9Dv7Oleu2RD9UhbgOT5EmRpeP
SqQbiGVTfjr76p8hCGpfq6LIhXvlVJWIiq0DH0gqSNC9U4mA0QXeYIbgsG0Rm9Qg868dY7eEy0mh
ll2ifXdQCtZqNYNBn5OiMLuCeUEKoCmJirf8mM1Ws6n0jjLWWqmpOXsaI3T5NfKXif/bbEMx4suY
oWuY4HZf6dLvQqouONJgWVmQdTcIt8AoWsf9D/36+6sYMQ2ZMYozaynXkVwzDZJIJhsDu+NF3pbG
xF+S1tF11oJzXtwRoSxfchH9rl2GbKKBEnX2f2KCS3sv/PESSdu4YVOSECD6Sw+S7PP0ZK3mPAfp
4QBdQjFDjE+8No8CD/l7kv0ALbqP4WpxvQQTRKexXyGGc/kdOlmOfRpXvIUtn8Dm93Mm7kpbkV+5
34W9L+u8yF3fk3ZDqO91Kpb33sbaJk50BtIpmnoz4+J6Voy1XusqGABwcRu3KOGkROT1hydh1PEe
3Mf6gd8Ewn4zuS9UvJ6SlkmmkwHQduPkOw50oIih0s458EKX3wzjVgZJCdG6fCqPeSRwxrhx9Oqa
RTG/Msm3uOqzxfHBy+InL0t915YqSYEGW02VN2f14IDMzTMsec3L89VUNZUk1j5mJ3P+QEdXFXRV
5WtkdeRNLaNg+C+nsrPkAkSG6LpD1+q7b8Qfzy870YdUnUlzlh/nHtDe3iOgcmD8zFF4Lr/XJrla
WhN3EUXdir54GfNKZ2x5V34ZxN5BMkFn3/HBvoECjC/4kh7ZXqAZsMb4qzTvhumx/VHg0SGF+dXD
7uGf9r2YHjh/u5dHA1YZeHo10WiSL6CVaMvxa1MAmsgzr7Ueiev/HtA+napsJlk6LHNOFsjAVFF8
L1sKYgvxGmeLcogThHQ6EKQOW32WIkIaqmL4HtGjbXnLDDrwV4wqS/ekx5WpTYgcKspq9Q5MY+Ob
kA5G/hW4sNfkrIZgcPze7i9owDwnwQTlzS10Iezpis/Ik0VOWm75gf9Mhi0OgGxFzrsRQdRyEGYa
rQq0Lg/Z2x2qqMA2h5CN2wFBvEc+L3ybV5BTQNqUDOvo2XR//EwiBakNpvKFrvHhvhV9jkZOXcrv
sQ0dSDALEXPxSwjhP1Fi5OOipIZsXqVJXxEwF1WS8tVUoqYzjSHtQostSbCzRuCxLHFJfWThnOYf
dMggiQUUTGIRHbks8A9YkhHN0I/YqXaKE+/sw2Y0G1qOpGPKGPOcl5Dc2MENbTXEbqSKg5DhL1yD
3AA/30NGXt0NFCOOTi/MNZpWyQD9liYo+RZQWlBq8G045sCIjmrOQSVeffYT3ddpL7ew/0jLBRbF
f18yycPBJ+5tAMTFryJmTQsdexyN9GnlWLxsYgzg+RIJpD27hmFkZeca+O9zawDUu8fBR6HEE9Ap
e/LDX8PpqG55nojekBQq2ucs82GIdZ16tGlk8TZOTM8NYcJzLHPjK3i2hm4ovhDHpVs5Z0kvX3/O
BqxaX7jGrUwfVw7P/p6jz1cRqAFUeyne6TFsse+UPWyzsC1lbd1cfO6Qrvb82CNt8wLHvdKh3GrB
6TSQJx7PQsbot/oP/oqUEGT3kVKRvw/BIJ7fK1zUVbvBfgPmRfJHeckrFDAY0lY0R1YebapeSFk4
vPWA077L62Pv9h93FdJ5WbsyAUCSg2yngTR8kYDvtgTQAThXmEhAN95yUNKMALC4/wTWeqKS1c1i
xqYKxvBGECCIowllnJM3Uj7pT8gDgp/BM0hNN8tGszccITsXUQjRI3cNflODo2+1dS3niqMYZmYq
JsekmePyyLpUFiWcW/IqJxHMKE9CVeL4rUpE2z+yjATqPDWfGGU3znJ/OTyFk8lEjo8EJqkyFK5z
Bz3hgdG2xA4NUv2L3zvHBu/JvU5eQtmWD8HaMlhWOGug2RruPmqc7CFn6E/6S67Onw+vDso7xvlw
Qn2m4DbX71lrxzpAqNVAsGk4dgcGc/gE1zEop72+AaooTrv0b1aMEA9Oh2dYB3j8E8NZ1UbUrLkA
6erBlZPEHicQd/bzS9sSKBV7X3QeqGsVC5B9RaT1Pgc8pZVrK5OMJhcTLvjoexg6ie3Fw2BnecB6
dvuC6VdvMIJS7ty8FyGH7ReDgQ8EeSugR8yWrxD53pkeA+b2Q3a7kOLGwxnBRIgk0WFOhGA1DEmY
xHG3BeIJU+/3wsoNaD/xyVUD00/z9wiPR+bEt71vvLs3vNA8qi+f9uRSgO2KmIzOxclDbJvPyy4G
bD3pibSwJYfXMWR3u1CC4+g24gu+eOlTnkw57/1t+IVxv3jp1ufM/bPp/KO6NQxGzk29UYGo3HY4
bPai38PYDP20HTRoDId5Q3zHJIZnY9uNk7THgHsLRXiBwF5hlG+P9s2lHBy3tT0G+7+4625t8bLo
KphrtmInM7NEeGn0Bew10AykhpwrtxNn89m4nIADeryOl8tLhCEqIZLAEHiPJiDTttJ59W60HpF+
E+Gk6qbF229cyjvmENeoO6iK/RLhlv/o7Rv9sAOmgiF5SiR2RQC3+/lGNgRmSXT3IZSxhUU3SdlR
B+FGeFaD2NTQb1QJPqJ4YgcK1zUqKbMS1Dgy+skpjXmslseKGrYQEwgrXxal6Er5IC3qa8LrVjqn
fkSuzGVj0hILlunS5nSQf1Kf4gpcUS0tWtO7SF7Sn8Ha5nCNHPlo9JWKyvQC+sOUGsvE8RnROqpZ
6I3lL0+nKCOP171o0pGNP3OjCttAH30GVzQr6fobGR/KACtlVYlgjCfG2KGMDhYYKWwiCkylLz/Y
48h+vtyjln36Ti0iIGfnB3qLUacLSUqwFR3eHSzZVEuCc7RMmkYRoNZ6T0DwnjoN8oVoTVKMdlvi
f6LSKiZsR6yy1n00wR3dV+KhU52hvie0OK79lGYtpPRkSIJqG5Ucp3t7fTecp+aKA/6yICb+oij1
/DANBf5whS8t+HmCZvrN3mIaYJxosf1k/YMYq1K+LpJfE7PhLPQxw1BHyXPDfgvR2TVEWhq18xLf
e0YC83GPsi7cSCnp9HfIwq+d9+xaOXzLImppHSAEprjfNjKiUrpk5zEKYXgyBcj9DG3SHAulccuk
OTt9ALFn1fnRRVJ9NWPAKitgVYQjW3fisb53PY2J5aBZaupGW/4wUgr2PJog6OiZtMB5TV++4Mbz
yB28PRaGl8SAC1hYiFU1JNCqDgHhc77SXBBmqb5bssWl8sPeMWw0EbiiRn26dKkjs8NLuLkdANm5
o4DjDEOrFQtSXjCgZKPGgMRK4G+cTl0i2h2HuD28cIDfhidXdhzmvSRnHNYGMP4srhHEZv0ec8GT
2LrD8h9Whsy+l8CoYj53rKcHCnmnrYCxDwiKw1pYth/L4r6KqvUAyC/Z/92dPI5b4KeAnQJIlJc7
sQQPOjFMp9TwiatV2ZQDLyrvUvNmS5SyI1FmbySWAkVoU+eTJbb8nn5H5VJGK7hNEi0QTKKayJpK
bFhh2cpXLQL0F+nSs5qKN9r+b97SzCwi5EOsFQ/M7HRLBfmGrfRB+KfxlcBZc/70d7XhQ3byEbJF
q1tYgLyap9A1QNZdwJLcopSFHokA5LMk80X5/0eHcxP5bScxBJZyJ4HVltMC2wWWA/zvKzqvKOFW
pFk42Fnz+TmYyo+EMSF2atuHCxi2+w3BbZafXcFufJwS4j42k1BXMfBiSZh/0v2YJP5FVcdHHat4
mmY/aR2FkXVTIybh4MUA5+WF+JEphH2tTf5wQ8N7qgezf6Wt8gPXhS3YIr01byXdKxBOs6vr5QDw
r1ZcQQSnOO670IcztMsXZS1VwUxHexU4LRsPysTtbg/2d0/qTgE1/zg+j6E1H7Cd5SSg1nCsLvz4
FcXLSxA8aXnJ6XlGdXVck5GAXi5FL16WCHWS8VWGMozXHNpi/d2Krgo1osFTgzSakdnmGDx3V94v
vxVDmlTeyfCyUAsRGO0sbIqph4qXIE2bII0/G1LTNdooxroX6Yhl3GoKEhOeV7u7nDtvU40r0e4r
zqlyiQ+IFjILj4imFQSOYpHOUjU4W+JHAmq1vBNvzpe0ttlxvqQQJWt2OZI8ToWNjgO436GdO7eG
Cp5iWZO84bNzaL4o3wyQT1bDj9dcoIm6Y6k2984mo9eYqqYanFfGwJ8utXFMTeZ50Lma6mAslzJ+
YjHuHvzMhyZ7nvOaM2G7BHyxeC68eOX2TpM3s+L5n40h2h13+q3J7c45bLD8f8HwXKD7h/x8uNE+
sTd1MaKYXcho4/i03+PseZk7xyyUi/lVk2Pn7DEFL9QAepZPht6Fo1q+iS6VSbc5XlHYiXewtGYj
21n/NXv8TjGZ4WmhxomkrlLd+Y2rntYOndaeGcOVPTOOq24i3pOaY1hYworX+PniRw9Y1c6mHlwh
5kclRWwChBlv6ZDPu45MQ51pq5G1ZzKF/+aotROu7u0dZki0C5b0bRT+y1GjzyIQw5B91pLN7JRA
VGhDjLyqRftCQwAXNnXF8e/Q9jdTP0FjgRq/a/s/Cl+D9hhEWy7zLEvo3I8+sFAtOPCyheyLK71e
fZYNIU8X+ZAYlXK4N1jLc5rvZv2OQamfP/IRS3/H9MNzotH5Cwc810MzBxsmoWaRy6ScIymIxj5D
YoioGMz423xmbvfy5gDWD/Sz1mpTMmdiHp5b0HkHOUzT1sVysz/mfOlD+lgHmYivtY4VSykIHH6H
IAWNuHsZrLMjTCbV39DfuhzhXewJvGqTP0esnk7m++PKKaFV0lAc2uZ6qO1Hxsh5JDox0aF+rMK7
DYYi/QQ6nz/m/hwYJs2ArpOwYwUbxQk47vf0PgHFPWlaic/1+WqqoXmJ36JKf22+a9c9mMWfq//M
u0/elVy5P1Zeewjh39mcSNCsP28QNn86AG8tgdQiy8VSUyFDo1Z3n5z2KxFVgwz72ikwf0jBj2qr
T04rr/MbX4zmJlW8YAMmmku0hngW7zubrGpUzxqz8d9oX45TMk4O7z11joQZq+KeBsK+8j6DV/hF
+RQAIpGQAF/IgYXRlWVdCPom+CuSHdhI0PV4vb5UfUn1Amcas9RXUZEvN03/wy/hwuXqvm5l5R6Z
MLkAmERLHjIR5rOf4M5VJoFS5r1vJ2G0m4zP7IdjK1JMX51lu7wzxQi3QdmuhuN0tU83uwlgE7A9
RjbloPuG6r0rxIkLEZxrlOprPvYevW4FEBlrS16Dzz1y3kWWr41jocHXyiRBO1UPHPfVwA6D0pke
8fPJx946J0iqLnbsoBUhz6kc/4CBH5LcFXnMtzleOLYyZc1pj57zRp/MlaQ96xey0EGMihTdWMCn
w+LOyIYXH0cQXrborYnKaXiqWlxcbx+iQDLK766Lxbz+xeof+96e6iGSx5JHQ/i0MFAFGmhhwuKx
kRRxLMIOq4j8sDiCsU7RHCeTNr7wP27SRr90/cNsXNqVR2T2XUjFT9YO+sfUbaYvLtC+aWF2eeRg
K7/HPD0/EuCzMUNMWRWBTBO7d7fAgC7sG2E67VicDz4DP/QbtuItBJ4fDre/MW4k9JEBwdJcOnwT
CD72vb2xXEPnrAoAS2/K+DJU3nxpZMaD20QNMVchdcSqZELJBpOHN7NELPR4WH4v43/MZKWL4cHP
75mh7Ksl9bfrubHU+WR0hRZk59nA1QvNvgmF2PkxVM50bJBIpWa/r49gFLG88ioJke8velTYSj+v
mojPjuxu7VQTTyjLQKKrGzG2qmG3nlVJUEabUBu5zlww65iCzU6p7Jcz784ai46rFxn44h7/WULF
un7DW8ywTsuz4co+sjlAe+NDdMu4Uzy4giuWnf29e50V1e/hKU1VvF2fPFEtJiW/ca4tIkIpvF3R
DTUieaSWXhAxzA91MULzQLKTe39qz+e5wL3dQXiMck9iiE2SMvyNKlJRbJUbdXhsHGuonNx+UA5N
rul+Wg9uMSJr99YBTiaFV9JnvsC5EWL9NE851lc5JY1e17Wq0gqz+BDsIsuYpkHONHUrTnTBLxiJ
HZUJJjd1zSucCQNMncGOx5rNcsrRCvNNUDB8TeTXo4da0samjTD9tObFACuuISWxSsXHMI2dfDSz
4JhDl4Ra9Zb0Br34KAm+jSvrCzXBVGL6DOI0+3jxKpVqAeBppJzlhygKJRbu9i5Wedes9iBE3Qm8
+GiWUFuANu8f2EJ4rPn05suHDYrRTx119VD9tHjqbUaLoWiuSLxLgrkBDpfitbVCbE2OsVSz+Q50
BzKl9hsunj5VyIonpTUQKE9Va0qHtTroOenoAWPGdFGGO+LOoZ1LoGP3eMAk6FjinDCuu+AT402P
9z/Jf58zvAnAUI6NtYKk4XLEoqrTKQ2PkjFw0DfWusMDZAom4xTvPpdoGidoR23bOLmCklwVni1K
Idpt62V9+LnJjCDHM4i/j7Sh3V3ltAk8hgeBj8qGGvSAlHlY/G0kGdID2o6Ml0JZoxzO4F5+LHrE
VvAdhRq7s7kgqF39XiwRbZDvYlFpgH1D5dmkQdloPFq1dUWws8zLFfxtYShOEyi2HVjtJldv6mdh
TzTf/nr9VtdKx4FV1cVXf/trzr+FZckPI/3xjRF6KHAr+E7jzL1exmIiDdME4CMXinOLWpypGRpm
CobnhrwtZ13FAsQw/uFlF/Qv1aVYY0pADLZq4b8vnNBXY/s2HK6eDHaM07vhM3f987PqcUpuBKy6
V+Hph1iHcLf6u5xoqhV1/P6Fh03fFIjOOcRcadZn1OsdWbQ4L508+c1DuhX5AmFBO5Y9kg6eUnHC
bzXlWVRGDftBEscJtNhZ8+o7s0SzhzyYS9atMxfAa5qr1M/5j8PLMLMvaKF0tHBf3heN0vsmfoH8
oHw04TWYx5xVbdaFhGD6ShexHWj9HeNp/OilnrcjnkXECOFE3SCtRCvgTTbY6Ysq4F+Rd4Nd2mPP
buHv626Cz/HqKo4cdcDdBTqUmP5as/g2FsCGETtt27PGjgbDcCz8iSQVJ1ppL9yNpkNdCGG0MTqj
3dDaYLsn/3ctfulfQIZwNrxR1hUmEmN36B+lIDgoYdYvmEZp7hiL5CjslE3MV/r3jtj5t/+hHgYe
df1TAEd9D/HmfyMTQLIZLbxL6gzufiFrnfi5ethnKfNQoFwRoFxIGo7t7PURU1Dnme5UcNuS3q6w
KrovfILKwfotOwxwhtxzEBE1EquyeYoDmA87XktTvNdY1ZMvlEd3Wu1PDo+BlQbpyMyKJWtB+sar
ApK0kxG6HpbbuudcZAYzvWIusU12BQCL+mjaAZPO8FNpvbz2LhTzIbnI9Q5SK7uYwqQyDtSxRa3V
2iNrkZfvb/p/jpnzWnM6VKYHiSICcs9rTlBCfr9k6tbLwKhmldkODSX9RtDEzoRkJQ+uCf1VlNVc
NLpj70QNsLqcxziErD+728OtXQ5MwGukkjFpx8mwyjLrwi2Hb0sTxGqQbU7bE9hJ4KjBz/zaYDYr
KWuyCKoUAAx6GJsjwI9DS45hwgvgvWeGV/2keOPLxBMmJcXPoNO2ItHp9eJ3TSygVQVrB2H8Lnfz
nHDWFtubmBypssNnIQVT8Bse+arQEKn6Tr91cWFxFNSlC2zYY3mWNgnhMNXI2NOwnlNFqfd93HGX
WBmAgZX1b+XeW14Xst3AKhtMgJ5GgWRhQUIAtRpPlENFPV0DZjgkfLYnTlqEmz5+LtlqQZ3oxA/N
AM0x4CYL/i2UOp9lX0Ki0baEXMWtey9Cqg/NwJilYgFt1tYnHePU3yp5PJ9Y6V57KfZ/IYFgzP4O
2m0KXBGAfTVeEz0NhGIYXbPjB6Yz3VIjaGxJg95BzqJxL+/lZXQZ4P6ggctqD++L9CcXuTJeJ9Ec
iFSEnsFVO9Tx3End8RhYTwdoyliSYUpd6tCwMcJonPB8JTYX9snCiEXb0oHIRyWgID8wkIDYyy3n
emiHkG+JOAqytAiJmu3Y7TOIfBcDxZAP04hrfrz6PP//KM+XmC6MwdY4x78n7Xevxl1mle6jhNZu
OkG8MD2DmbKZRclRIbbI2mEVLJ2lChlX5GivED14WK3+ZR3eoaLpbuo26wVVnktFiNAVzbQyFs0F
QSHEGKv/5Ruo94PytJZ1HVeN1UtQxl+/R/XloIgFvhPKBk0YlWKwx8jen2h3bx3bg2tRxXiH+Grz
dw+sJd7NKthdlvlbJg9SXeZxazKRB5zUZQVe5jrFl1egDCfHqPgQ76C6H3rhDnV/r0LfKd4NWqd8
OJgyoNFkTICSpSLeldKVvZW3mmMCXMlKoofz2+xmgcWqEPSyX2SPIZ+ngZva9r2elZ0tspZ5ugB9
WEjFMb9H+kZYwqpbTrQF5ptMw4+5I/dCJR1/qOgun24kndI+EvxrahE7enbjj7u3+MI4s3r6S+FG
WHjQgOPpzabvZ7HgiED3XuL5Qp16xwMi+UyL5Gu6nC3+Bn/dS5sj03lNghIO0o4qLB1f0EkqfIO0
CS1+VawTifS3ZaxXK0UwDgAt2jfz++7r/DHUO4MLk2b7IARjvAh2Z6A6oRO3TNRowloht0nyHjrY
V7Ro9xW5o0dgYNM6/RWizmM13Fz+iEn74+uNfWV8yqCFpw8D1f2lxmnixqHxPOPBP9kK30N1L3hc
d1lb/8w5R6j5pWRVIru5D6Q+QT7GDQR7YgOpTNX4Gmo7lltOMZRJP1OQxlMZLcmHar949D8NQbPn
/qWXohFyTQnSjiJZtlaPmi9G2H0LCVjcIwZpYYHs/ouHhU7nLVMfG4E2MMVAdEJu7bXJxz/ZVsSW
QICbvEpACREQ2+hsyRUTNcUD1T4/+1+xS2qV7R7mc3jpQy1rnWA2AmWHsjk+KlBP679WALX0w5K7
U+rOYTPE8UMkxQDjQHN7oKeLuEIcmipTvSDx4Uspx2x0nl60fIIFYKG+HAIN/ddUrxrTXpkAqZhO
FXjIc+Ot302/VINlAOI/w7N2qtaKAfpMdH1gboZtOtUUswK6IYZdP7HleQyW85PMUqr32+11EGEY
6zqp6D7DjYtXF0LBwJ5KWSF4+DJHlm28kXelEtaBKrWKyA89KHbpNUQOZwl0I17MzvXh92CmjnnL
nfyTqT4f3NrI5cRKv+70FiAp653cza0CsX0d55DeuV7N4+jsUzwLO2LW4zLW335XznSI8eyG8rpx
uULWjo144oOz5tEZpsBMBYer6o20iGAbW5o1vkrNIIAPhUTgKSSmYk0P7SoFL7mMG6zxxEskfqc4
VkKKj2gd0k0+rG47UmVe0bAWNmnj76FW3CFkQ79r+OIYQ2DceULGh4PnEGTwDvQaNBq/OUFYcK+X
AMX5JR8gA+qamqsd/NGP5V45/7GmNalvsI7JbEBJqgF3oJH8XHtX4WjbiUH3ksSIgx+EIzG3DeBA
2etCkP6P7woBFEttkwjiL54piDGuShZQgbqLmSpJtUB9+JiUxHEVAYvqwZorc65sBvJIjDIkSwqc
c7J1O8ScoUa8KuqoDomJo4VgKDWZ0RHRvAYC3Et6bOb0iM+KydJBs3ESP+J13E0RA8v4IKfRBrcj
6Tc3Qi24C6mLzGT0S/kCBMs5FCEAjDGTVmXoZ+cuQSXnKAT6WEPeJnS7ktymFc6RuF1zFJilV+jB
cGX3VOii6oowmKLU8Xa7sXqRfakkCCX40BQsVlFNcUOp2HBalDk+66wq4M4eGB2/4B0jwZx4LwS/
oL8qmnYk9BxrRiuBgJJtDBTBy8Hj2Gw1Kfyf46wHSNXbWEzolGiuX7wfKiYy2v/Zz3z/RNXlHAqb
Jq0NYX331D5gB+JBAjzl+DIi0HxBer4w1ADg3Il1xHQxoSqiaukMwf+OQ5c7CbvJ1cplKQRnZPtg
R4YDjtdLkCZTNSCGaD5TeAgJkmU3VbUMrrqrMk5Cg9hKDxk/ujBfYux7w1oVownPaj1OpFs+San+
2utuQaqoFeLvQXUVwMJXCFekrFeNiWnEwZzQ0+y1zEghF9JNd7N0Fk9qhe+ab2Ar/OY0Qr2gCfNo
UjyJtx2pIuJCQYmbICXJw+k3zSFVEaMDyRPsxDrl4ltKicAio98Y9eX60VVI4SLI3FSKVzOUaxiX
fmidHEQORwTq8Z7wnsqzDwuU3mBYENZWBygAhetWeHDFjmEs8iUbOZO+L2YdbJWQkQZN3lymktRV
NXqDuQyMZyDN3I92EZpQQmtSVRqvlmRRpIULXXocyUlbHx9CakmYsOebCnvGML84EsiEr+cxLNlB
beY/L2bQcfehKE1t2Qh1W0xUPqcu7EyZr+DiEixPfsgpE8cU/bOorLmZpncx8x15Aq3VPjt/+/oc
o7yrTe60p/wQXTgMXlZ4tnbWdcyxxcQ2d80F3bPjMLHEdAYWMQmVXCQgyhsW8gKA+6mesoMq56KT
QO0KJchV97k7454+IkZBr3U8ztHN48vC7PAxfwzGb2HrBv1haryvdNKO5akn0H8qQCj8Q6XCtVH6
zMJ5UYcTK8XNPHxfHCwnvAx6PFVuAm7KdGl8u9RDhTFpoDPGlnGgkOsr8RcrXfuCdBd02dsDHjYo
6AydpaHMR9NxTjM02ENiRKRFoNsTQflxht+UEHfzlhSF3lPAWBJFnUzCVT8yrvnh40CVOdnhQNhj
zf5TfMFSdCEYYAduDZC64wwnhNfqEv0ExnJlqhj54h17e2GdjmLR78ajrzYWWJ7D22/PMGDISlNd
zxZkpy5BhugrvMq0qgdqxA83S8PCqNBMyN9X+ZIHeDCkPyU+mcJjBxyiH73wgLNQj0hEmrOVDQbS
9GAzdQ8pT2MrU0o1EL9+paZY5ak9DAtZyENF4JFpLDfhZ5iTaDi7qchnKneO4d215CxQU4Ktqz83
pWDgy0fWmpBYmqCUvyYleyEp95a54g8tA058JBZEEbhSCHsXdQS3bXEgWPeRq9EFTurviQ9tJvAL
p1ruVdvBMwq5RwNJ3KGfK2w7oeozqoBB59J16C8ZFtwurzwrvT9HrL+4dCzjhyF8X9OCBmG+SOhl
FIZZur9UQ9TFEItYPH2C+he28KUMV6YteKmTAPzH5h7HsebbHaVEJa5YbpcZydX5LHZrjUCiInxw
KTxnZQv2KGPifYhP9Xq+dbCKgJrKfkadwuCoz8rTWhpTIgBLhDcuWJWESp5ryfqO1TRwbZGX128q
q3uKZKNQZZatj+AmIAnywvnf5a59MwUHjf4OcRYZTs2ErL2VohpO0HPspJ3ZhjquYzkhBwKZX4TL
xJzVpcvJzAdZPhwqkLhaOj7sK55+Kiv2dNYAokcTZGZlCi693yphrNRE8kSAlK0yMFgscztsOHpR
uZ4WCKsl8wy/qm1hFYlo1YY9euu2bCzDCFIOCIDfRMd27dpuj4kEpiyAV3iBHbMMd9OQ0tjoKUoM
N1mvWAdxRjF+7L4Qzh1z+2pGbtW7doIfd7un3pO6oRaBur4Ngi6+wAYxTbPA94CPo5XVvujGOhTm
bNC6oqb/w4svakNx684bU3QKYqBnI0PrzYIMBuHy+y3VZ0YHRqS1BoNE6gzAHugI7xxTi0U3q9lx
sWk7ha3uMr3MCJC806dkaOOSZpqYz21VVhzoGQ4XcwTYakkNxcYt0PiSsxRqsz3SH4txHasLzSyq
dTscDYV1jmXdrPeoarj5GGrHhEeu3/FNg58wMjtMEbl0YuMxd1mKao+shyZoBz4oxtvrxfQmET8M
W01Mh5etXOcWtB/1I/GEGrzGErnnqC62OuCAZL0Uv/qT+q6SzVN3nHETiM0XBwDMhKu2S+RMo/HR
I5/0DE6JAJPRrx/DhV/n5z4t5CKzapHv1UjdUStpaYGLApyY6RLtT+Ivs+6SZaVaHXy9l+/egZV3
cB766rNRK/uyHJOdrF3CloD6lHpROfk+S3OIhklj5kTh5l+uu0T0e9pPc0yMAuT7URzqxKVYNp5O
P6iV2o45V9BKjqg9abCmjjaw0GbQ96+SsP8qNmeTJMLqFRP+ogdu4vLqZV73ba9OA/9J/Uq8HSs3
NXH0/anW4EmPoFUgqLjgoX6Rezb5qoaepAGf0eFpvkKcfK4FMLairweM43jQGGtXKaj5H3D6+VrB
1WdPe/Eov/6bjCKhPuzm122l2fWP1IZG7cNzVvMnQV0BcCFfRns5tfEtnw4Puxj3BnMOVMvuAsKD
u9qj5T1bqVKGF2FEZcewA0aH4sKBPsucJpqv+MZRT66/xaXG0db7O6ZzzAEtnM3XJElXMiYQ04SD
GSjU6ZCbHcl1eBTq4e9+3cVRTFwUvHm0RjHb/6ZQwcmA3+qzlnsNYVCe1y0sXUQLz6wUhESqO7v/
0moehq36EOA2tKlrmmghDYErhgJwqKYKX6xgI3iiAah3hxgIUCiWpquGpsFyR4HZhUWVd+8v3bP9
rAY4fpOrHxBwb2873WSdMZCRVN4sBu/S7Qsibg8hWQTIoiwbXtVplU32YaRasWQp0UhAyWr4Cr8f
PztLZ6jY7ONZuO4u3FLkrOHEqPL8jSnmhdq2rfFFTdjLjq54HP/nsFjjby1r7U4MBPjsYGyjrlwm
UoK2ldg8N8Xcuv7vn4xdO+5DpxpKtdvoakhleGOlTIjPH0/rvj92nLMBsoIAy5wZE7A109Y3Ta6d
oByUhWki4pyJ0zgjIqMCLM9QvV18RkhLsVuzMgwEc/JFkWaupV/0Zp3+5dYrc5XvmDz2CrixWx2d
7AdFF/hJR3Hb+1IaeXhY5F3/N/B4KTIXolbD7KRP8ziUmopFKY7lLSxEvtqJKE+l5aFE7KpdR5pW
gSJ7MYswBp+bj/EeIIPEiKC/QHcQyoW4XuXKm6QK7g0B0FxkBakX2WB0tO4bjXWvXCnrj2xQA7qU
EISv7XUpwrGRSo9hV5DfWqyF7IAkeKHeoCyT0+MzfZ0kM0j4NXguiVjriNk8zIrvw54YRTP0tqi5
vPZxCcX5sPuEOiYv3H1qqIiZd9xh51IqBice17JKl7/slpnCyuyO3geP7T1RuwVUXrDpBCQiqzhG
l9scNZ8YDgXWyt9fDxGBIF3fN6RbwRSuI13+NDQxVs9wYBTleo/ni0kFMwfuib8KN49fd0xFWbfy
Kdkc2F8EnxbwNnt0aHMwrrj0ewWxxKvSPChyCc2zR5fTBmcPH4z+LVeQAW8vo9WWtfkLQssHv/7s
4GDM3lhTdinMfSxFJWiVfZ7Ct9Zxr52cr+EVr/yddzWvWa48G5ktvN3hTsgvo6KADsqS5wfH+tuR
vj3xyTDLl1QWhD+5nzRzfUj0PpKgzBkutVCsLmjvbUSNQS6M5voTUJDZzQrpaUOEFe+s9kh34E0i
LUrZIL+3kiICsVM4/6T5iNdQhAp1EybUiLDPmTfyutXYBzBNgxSzW2Z0VY6SFtXmixymznbU4sZ8
A8hACZp4m3TOHgOV4J84vvlVi2p7W26LDrs7PdHDrZ28e2MofBLzHmW1Kw+grlkeeC/n34hHqQp8
8eiLX96RVFN+nx/J1gz1eLiqz9qVNKfqdszYZCNtAKPla9+n8qNyO4KfXVLeOMqkALTkRbJF8mz9
pRDVZM9kXZnVhWggD5lOxN+pjZJG4DWAhsP/cT22VLy2lSA+uIvsVK/BBo3hATx3PC41Pzqr5lAo
/AaKBwuzIzpwl63L1meEbPnkgCC/FccQprEPYuAz3zbYp7uojr8hlF7wY6SXO1rLkRqoi00tJUqT
aoKZdDLGT02uf9O5kbQDPinC5WlSOZmyBjvdy8QT3mH6YwNm/U5/AhgHDSA+gzUl48OaZbLsDVk0
OCzEuCOPu+iN5U82QQuCgk4rLBV4Umb+rr060Ey/KmiffulnHl9GnxEfVBcZhE2nBtPz9mj0TjfE
+3C/goyPP72+FZ4HMXZ41/3lfFVVRpbve5JRcb3NPP+e5KHCzZCoWUFiSwFiJNRNfbCVhDBVR8m8
Ekn06EQoEgYyoLAKTGHnzhbiYUzGpmLIXPa4KI/MUb7CsEKHbWzb+0Okvw00ITTleZ+ft5yOC6To
WtSYT0F1Tqhar7awq/9g/SMMp991ZA1xb03wB4CqE+mlf2DB9vqcp6gkSjQDXDQW0l595y3gnHa/
ZohJWpmT8ca8FStSv1Ml0orWN/XGuzU+O0saBEq64ANO4XUkj1Obhk1JYTG8pA+WXmaAtJ74MBiD
2ux1DW5wCLHcGKks0Ta/kZMMFvql6fsbusvWAZJfZNg3xwETYS66XJ78+ICsRhv1OxhlPw9cKNuN
z2qYjGCC5cf9Pd9556SGA+InUaxewoIRW86fQ5j1af4CLlcdJJnpfD3yW2CInBKEIEB6kxd/Xvxd
LoYEZoGOCtLCLtvNivZwfVRbkQeh5Llhel9ShJVYPJJ9uZ4m/62+cOfYT74UpM4STMcrivwsmgjI
x0OeA2onvw4zwBjp6GcneuG68rvKAKsugzphptCrXcux43HSdgOkfe0KU50dvlaEgzo9fX4sLPUS
JKKstdSCf+0W0fO2aXlIKWaGGyZdFJGLATma0sqJlKa5rrvO01hRhTijCddTjoZwosq1W7GZRCeH
JV5UIQ3/HurHccB0H9FVyA34Pw8CeogirrL9j0waN6eRp5tRzRg3uF0+eyPNMlSxUn2cqzbuQBZl
TIpkvCBycMia96jjSLiZAKST9c1W0HPtHp5gvCFmu4SDtV9wKG+uGJ36p4XcWz/WmbDWQCRtIh4p
wKZM0hV4wlz2kxufN+tskIbnMULXe01yosgiBkwd4jn7H36seAmGAJtiTLqIU85q9j2eCRGoH+EH
aGlmEJuFGrxqb5jsgnfdPwR6irMM6ahYPrLmjjhhWrOh1fe00/2i8FDtDv3MyIXiXvjUTaK2JO5B
UbnlWwKuOnKQZFuH1FHd00aJ8NaY0v+f1Sz/Qr+WRMk0GrOUFqgsNVR+VSVz7v9K1OnaRpwKgHrS
vPVdzZ8Tm5k+89RqiEd7IiNyXfO4lGrFvnRWaEOhPHKVGK7993SjKty6pSWX/gu8j2ZbrBuWEIz2
VdGK7/HNd3aJuz0ywVQ4plPW0Dc+2YV2n2MECweextf7kqXrWa5djb6ilVTFWGV4TDNx/O+qgnwP
Z4w7tjRF6DbE/TvOjy8zNL0/8pXQsBWYesdObvfgvZSEDF69MNBs60NqhsO83zwjZ6G/wFUiAeQ4
AzAU4E7N/jH0RMrbqQMA8CENeuxn/vB0xOKvgbZmJBieWZwinhoS76Att5336oQi8MP6paIGPbva
xUAx3SG7azD3Z2qohv6uOe682oh4dobDXqrsQr97ZyCBdlt6iaXtbdNSADXmdYbe4M2VuyWPgtUP
2OXRjZaivALlESyMJy6uiK/9cz4H6JMJ20tLfeQQ1hHn1VSsXUWb7yFb8XutZA509t3T2LazDRZV
yMri9ttYkB3X6JUp0B1p8RjaQsX6smGvRZ2NQop7jSndO8cAHdZLLj6aoaOHdEJ9dkU1/ix2wQ3U
hKKUlvRuURntMTEPxT3lDuqPUews4y0cRIhi3b0CnmV2CCfD+wUaGpBitEZbQYGSqDKo2ubSairD
v7ENsXbHpkV22XXguE/HMjfUtB67hXR3DHY5heLwBL+yxywJuKgb32mDGllg7kICjfPnxMY6qIdT
+gSMmhF6vcx7JrevgTEOMzDMWQioLug6q0W6Kq0ct2TXCnjhKD5sJTp+XhFyDpiRaWrTUq6X2UxT
XO75DTnWTN0xRcm9L7mAjXFgHSKPAiMEzgBDOkGpRnwea+TG061Kkj8PxeHZmNuC1tT9seGdujow
nsTwMDhEzbNa24CRh+xEy43eDdob/lgkRHLu9Y4Z/1NtTKGX1M3UDzyIGEmvBLcDtqtyBi1HVTPJ
lWa0esD5V7Vit/8XKXPgCofcXp65TqfAPR3Y1aWIOc/9gQBTXrwY6EKSsXhfs8yuSa4Z0nAfDliH
YEIj0E0oAj9FO98nNf3yt9bLtKg88cYJ8eF9CoYRkzpbgq88cE0WGQ+X9756SoFnQ1pnqrYK4bQk
HSiHaj6mMsoLnWwyK05bAAjNu2LnZtf3CwUJBAXC+8tJLG68LX7VJAVw463rEIsxaurRNG3lHvhh
JaACROV5+q8WYw+cClEKhMBAeBkxhVgD4GIXQiH6YCyQyjmyfz3xQ3SEmsRxQDIKYEOP5IcfC40R
6iqcWAfN+NGcx+E5yUleUa1dxCgPCk6WO9WPTeod1dAsYzuPWzSb2l7pgQ2RRQOuxW81bQ7aFhFc
0/9cgJGCgQ7Y5/c8acivejwSpYPYMHLrwkWRt9m53a6eacOOG4pR8VJD5NNa+5gE/7u81echiHPZ
QYQnEzbSzufeShtCDuYmsJrKzerdTu8cgISuOBiBCtmO0S5B5//eIWRJ+0nwpIZPwWn4XkjnVTZD
x4qt+J9x2ogm/sbQt8lN92QZwtM3bkFUpNaY41eRSUgS7TBsOzRu+U55kmzO+c77s66EsIxMsVq3
nzk65t6uHZSE9+YzD6LYJiHuKW06Fa7VF3uouJ7pD6/xMGk/yrfDA5Eywn8Mv/LLU79BaXGDPZ6m
IXwX+aCxCrbuyiMhi/TysBEx77CLOWKGeiSFaXRpHojHLR7waZOWJPEWc3wr9t59qHxMYSGBc/6s
UEthEcgyFpWuWeUWnEemA8MfK0bKg6Wx89TWOqpRBdwdsoWFOvx9S0JPckePvB+fjn7rBFOr2JEK
hxs0md8tmiPCcn4uNsGakWmA0VJ1KXLp2Bnyp2ymyuzdE4YkdsIgjx6uIU5pbxyHK84vftuet7tn
23/WKWkWDCAAhjTnRWFqy/hkGrTHCAEMgYikv+gybyHpKjGyhB+ypfG+r7LNvrWXV0NZ/+y4BOKP
gEBJ/UKHj/kdaeyd8NUkIPNoqMmcnKUD5KnUJLRCbk27WYWHc0VQqKSs4FgRNBpdoGoAZ5IMLjCF
Q7h5OwkSuhAUIN2VdJFABghjrh6iVIK/bJXBSmBvUNORNVsViVdwPwy1eDZ0mn7k9zVNAnh7YMDN
93A2nzmg1KVumM49Cg83u26Zmf7DlzPgPZrEuBSlmXhr8WsI7hmmBXvAypo/Rx8CVW9HUAW4I0XA
0cVX0114DpODgLvQM8qF/gXFt4XiIVWZUPekOPBlqYy/taz2rxz/s0RzcErTBBU+nTALNvPdtBv/
GZWMAAjTOp2TFSFowWuCPzhWWPZIziZEr3uN0RhYNhcIEhWnlmsdnb6hdVrXpJmQB3VgNKcZGljQ
sghfXVSJGHxWFzel9nlqdLVF+omHSMFp5eB1X8jABsbNc5gaXnakUJP2gSV8AI9ASJIY6tUMVc4T
DXExVxtCLIFcx8gjBXGpj7Yenes3KgBubkjXW47afIbyt78fejz1QvxZZxQylDsT9eb4LaqsJ2Af
VLUK5ACUTc2qvM2+w5t8rABbtIovc63veFXECyL5yM8up9V8HTueab0W6ZHH0LSmqF00DNCTs+Qc
A/AzieBOXO/J2CIy4vv/GARbizkOAewpytAGmVB8fedwdCRlKfgV4e0ahru0ZtzFet4Bfz1vv30j
NXC6/Bh7lFguKqKKcsi7Oa9buQ51gWtjfP182z/s61tcHQUoZCdT72KqxFUAztewORlg1/Xj1o8c
o3pN8LcIrQEmntQm6eV2lPPBHP/rNDLHMMuODKQb3W73Enz4YoYhNpn69RsAQpo7RIjGUBokNKMZ
jR951eWzyhe9lQiS7gMJUUEyUfUE1gDNvZiExkiU+iB4XWnAGonSHyzY6xSn/g7KPZJXz3AbdMkL
eQVcGz0Omfw4tejsEp/efwTpXP7nZDsnAqxolNWmCVTzvw/i9sPsfxhzO9OgqA16uMQcgfjl7XJS
lkpIyOqaxWrWcqAhTTwdQS7Hp9HlUbnhoaA3/l8pc0LSnc/k3Tp7HrQZvTUwTywwagu0QErXVdxp
3R6IY0kMoRMYlbAyFpc1lrQmxxuyu3UxQuXCu4bmeozaNpxNlGuMyH03oaYu88pCoA7/F4uLNQcL
hvdWYiWTSQbeUCHD1WdZ3mwrk4qrrOus5Hvx8nMY0OVcwnBqJq1AUzPnLUMNt/j7815I1YxUZI2T
OKXKexNCBI6wbj7LHiaCVPOo5xtq4sTVrD3YYa6IuBJdmhBIilMjdXd6CrJcJ7/QzrowGACs28f3
l2vmriGIUFPO80E7fz43orLA5pLjh9+M866zvYIJI4n6b7qNpiDDp3UOq+v4QMv6MB1CrP7jiWb2
ZaXWOV96lnArE+TAevQRXDwA6q+2bVSz0x+WGai+H9QkG6ntFpCh83YkF7jyvKB4BmvkQ5myjS+/
UlbZbDS1xCgiAXgKZYIt3ykpjLf3oV1qvCyPJ87r0R2Ld70uGjYnZB9FuykPjVi98idFMong4Bsc
sEHAdaz6A9Lb6eb4cuJB8rpdHjIbzXfTEZzFxn8o1ztufhbkp1tvs3HS/+HWal8Ur/et2YOwikiP
NGDd0xSE8G2YiXlcK/+8+4Dq2bo5sImV+WtOzlcZ8e8cwkF2vYbRmZkNjPUFLTAuArV9zYJaSJW4
IdyoSk+MtoQHEGxPqHKk4bZHAr+xfE3XM6VfgAH/05ju036JO6mkAn5v7husAnn5kM4loZbBPzAE
DctIKoweU19au0XK34wpnBYgmI8MguGEzQ0CB23sjflx7D6j1FHrpOYLLi5Q1nh//tScBJGeKdsG
kkbJ3CSQ/rpOPWEygej5/xFR4M2pDDbCrzt5cIsEPGuVeazl6YY/xpbyAB7/pYKNXN5Hrk5oSAmo
NUJNq/vn0cIrfgBc4twmsptgP84jakv8tXvjHiup4Lw6P5KmBoJcRZwQ5e31GYEaUS7/o0E5u/c/
KKMUn7FdEffJ+HjH3d92BL+Wd7GuKY6/MrG+WlzvI2oYn5z8r11fPJymbhlDw2c8ekIGLG7d2Y2d
0VfUCaGQ8K8ifEYC3Pny9yEpnMIgVw79MB062XbGllcJPRznctZZYt3xIRHc1zkgFUkdfS1kHdB1
84fLNFu7dQ7gcb5XmPmUViWOr2w68dOVKCVaRRms1xAcJpTo4KIwfK0m1Sq/L5voKx5uDcf+DfYU
Q4COegjf8+jFAax1P5a25W0HZEPjZuduzs3tf8UU3O9UHyvePz05jAWZDxV4Wx6qn059r3jUPJ47
bq1/l7YZkVYmoxflwj/is4P6ZNRZdlgVcRhLk0bGoCQr1ynyYpP59qXlOiiYD/vPwAC/RGzF4CXt
FHrdQOYT/tsxsTBV/SW8NUPkko1j4i5xv4RsHTIYHHEsCuJOwgfksswy/dA1aSOu/tIiAr9Bqbs9
GrRdS+ehxvHsBNW0pmvp/rPmJZiNs2MUWFqEw9iBUx/HNbzolEBMVis9l4b51Ya3JjA+s0xVmWIn
fXkjfar0ZVtRTtZoRkFoADzm7Ef3cDZLGDJWhtC1DEDofQIxu4UhJEaCH4IFF2KuSbFQPQ3VLvA4
C9Yy8T7aqhwHu72h1saaTYv2nvxA87q7xRYzS9SeZXeHknkWgV2oVlX+E1oF1G4Fih2rV7znWckq
dJCWz84kkwIwUnk5xcamyk8qNuji4NlkrnRAAQdjKXBOqd1353zkBj5/tgqFmm/M26hhkljwuJBX
qZ3QJrD1vZzK8qGCH0dvk66Hx9XQCk18Fn5YOrB5hfH2f1bPV+S2Wy/Z4tsvEdyzQba/rRyQBTp2
7tMhuwDvPLSvfQ5oPXiQ0x9zfz2j4I/nusIgqAu6BU8sk+TfN2Wf46qaa/+6jYPqio7iRj+zKPwW
Xx85PHI4WS9XQurjODIncleLCV80kH1tY0rw3axamR1smknEQkmq8uc92qGFlAaZrWw24F0q7kv/
qo2HkQJ9HrvlgKmYl1c3KdScbFCXPQjyvYvIaaHmuPkN3o2bbTjiuUNAKm8FVXRidvGzqTBesLbb
KVIctOhoSX3OsFpdO/K5YunyeRhioJRnpuYal7FeAcKJbca0DxIejOek67X/6g7lQXZqt7IwOdex
v5R7sS5fL8kZeWyafGpbv/bqZUFBceWMzCYqYtEbIljgp9ghB7Xx560huwNHFo0CiWFcQRyQPYRu
86hiOoFQEHnsaUbNK/ycX1MseI20A4X/pzYvoxkuI00tXSXDVKKr4YMJn+bOGRgN1ZV66JMtDclb
oRP7Xqn6ayx6gmKyAX3bC7FZKnXW+2HunvYf2lHekNFXnz1JvL4D98djpZsuykW64X8QVHZiZnxb
e8x/gbpkj9XSQua1w5hDe30m9xMXWUJd9r8+401R0mG2LZkDcsNtMadHFi9rlGPKuBYmczVALxya
41fnEasqPEPBEwp8Ei9nYw3pTTGABd+dVjKUQEPUvTpYKc4b4lEbkUzETjo+ohGjGPPsnKuWnyYJ
m9s0vL3Nf5Tx7vEBxd6u5gF5Hx1z3LKviU4H9yK9uI34KrQgB6ZmLWY/S5lyHJM83XDPE3YFu8+6
G3LlwB5HoBOZVrmVosFSZZ3MD1ZP7ykR2M4vhMQxlfUeJwq3Bzy0OkmrVp9N9mshJW2gaDHXVT+O
LCtlUTexGOlAMQjezsSiSz+ClRTIypJIHJt34FkDjf4iQCTNNcpuO8/AmA5mU3kWHx7TixzVzq0V
xGHk/ZWACnpL2Fz+CDKraFBLdBjhNyk8FDdloHvbJPINLw/TGAyarFksug7EnvHYp6pqKT92fwNS
mC0cXTROH+zR7XEl0HD4SpZ8HOz7KPVAZKlIjUmJyWgFvBprrInbwInu0Z7QKKOi4pTTqTaF+Nbt
SEprvyx+Z/qYRw1ReMFw8xWonPloECAx+LMjMaL9ENTOXAo4ceEuSeYFCv714oazjvNYVTgrMOIv
0jSiyQJ1fkSGMlDaQ95Tj+j1UaeWV/0Wd58qDtDM80NRMSoB6zsdUZmO4Jw7LbQvWcb8IDzmcGH8
MJVRd4HAcoIl99IuNs74T4k8Y/klg669ofH9HZD279Sdyj8sn9NfQNiEKYg+GRrqW1aI5z8zeUuq
W20B+NgvaCAc0+G3xa2UIeJeT+g0OobqQks0B5bXAjaIb3y1PGy7vJ6fGa6cZ5yCN4R5TLrmK55U
zrCYytu/shNfNmW6earNPEuEgTRFlN4m2qlgK1TJHIlou9rpAl322JwEdBIXlxTDO76zh8mJGqLd
C6Ak35NhLuN/sCYJBpN5tdcxsXpY9MQlw/jw85IHqMmPl0wICSxMy9PcWbAx1Axn4aPFob5FufjW
8oq1BypqBolBhLS6aDPZ16bLL3jVRepE3unR6/WX76Cnd2U8zAD85HvJafxG2WHYFVQ9gtPWDLeu
ubwzTt4+XUUnNeq14EmHz6u7jZv2leKzojuqf/NvVjvA2sN5+Kv3zJIxIzexG4542H0euxE7cQ9C
xUtSoO343oKLGhSQEOCWWiHI4VHk7Lnz7PG/SGVDSxCVry19km85koLKAb3WIsGg9yE3sVkFZeJW
ynY6HPfaZ/Dz0GEI2Fsaq+YipxtXRyy0AcCIO9i7z1Jf+DcEumeLpRGLXMNYqK4XBAlT0oN1rX3c
GDv9c1HugAAHk9T5kaPQCbAJADpcostrUkyyQdgj5PvDUeENyFD4rucJmREuCVnZuFrudNg6kwZK
xx0F+Pvkozpw9Kf7xo7iyfB4O+aHjsCxnCy7nErn//taoTXu/bX2xg+Q6gOR/AWrYYDsuQVxPhqF
03/1FmEpgeQmLdd72Id8Fg9+8IXNZB6N/UTBk1i7IOWY/xhBbqOiWZwk3dTP3sRMiFQEjE6ue9NX
g+Tj855IX3ct50bwruzRu1zGL/Qovp3tl/Ncpuj2+cXPelwqq0CijnGB/kBufHWkcosVJJJ3NjY9
91yxGnrdqEsYxbdNo47nDnb0DHGoGNvhFOJOr/jA75CkpZ0kiMW1nOm8QmRwgBmGAEZWD7sTivDs
ZFsUgJe+Ub1KVezHL/ZaK7wN8/g6pjQSksShG5+SG04XMk7b1yVTHFTHc2we8UaXxrN4T+KAc2AP
gZOA1bFWw/ZApS9TF5cJIteovtNgNC0vxS0Ghlgw7ESEsUDluCqDQCr3RkO9Yhl5driBK6mgqWwF
eNkQ9DZHlcxyZSRssDitk3AlFbCz2I9BdE78ZA+ieZECDVMMjz9pPpTuYm9I5BFBnpAcnHfgO9Q6
qdpKZEI1qx8Lhp/Rrf88VXCmMMV/Z4BXNNEfu/ssFYjvlOC/dTSXLepgVK9Mr1sf0KL+SX7i8vso
bSkBEivvmHWhfVRWJnYDpPs7avO6uTkJse1+PVZB4kYZuZqxqLcDgzUeMw57V1SF85J7F29OXF6H
Vc3K/gIeuDYmEjXcvhsQxwaVfDiGkQo4QFY5gF7sSenpbIT39qRITNykCa7/Ht/hlpvZX53RJ5nB
WDMZjq8wwhljc1+7K9kfQhxW5NGGvnje8ttN/a8fuTwfc/NkPJ4oDqw5UjnxbLKr+F1EKQFZYnNU
ZQxwtVI01e7BhZ07I4qtpc+TLjFYw1gH8WoucCJjnn4oLW7psB023Rd0Eijptlzw+dw8wSunTAmu
V/atjVQTnaxpP2jaSvwGDczVyZcEc0ZplFSIL53fmTn5iOTeOrhp4UxXmqWJFGNxX1eHMA4CQc6U
hdt1jItcUUEUklJCoaEt2t376yb2rAHl17ZcXLZEUvuFF9CYLoV1sxyn9qKtRYFJ5dcy4/XZ1Hsy
xk7w8F5uLCuVtv7cFPGZi+N30qBRajT7rDIiJSUc+lIxHQPK6gfySd29Vm2fK9XIjoi2vgi2MbTV
Hphex+NZuyu33TI07NPwnd6zSsm29OIk/8OZ0chXg9ps2wkLLmjAsmXqa7mLXXz1Z7lx7POcdnRd
hBGOPwwP5TbSQQM7aA4yLCuBG1ST4yUZxVl0Lkvpp+d8+JkO8QTGMLA6QUA1NVjB2YVTm4AcK+2l
OXwfaltjUhGxao5yJIv9oQWd2fa3WKZyquMnaAdt2+zH/aFxYR8PoTYOB7dV/SCi/9xDJsTTUlxL
YFNO82U9gTB7pAL7CS2gOyT9fvmutnuBxw6XZSuSsTev6OpE0nr5dPuzeQWjAUodI+6l6umq/jam
WHlL8/4S2SI6qf76dQFM/5+A2fVkdOHsmAZvpGZCCt3s2E9wKglr2LTdizkPFuEBAYSGFiw7peRV
7qt/C2cKt8ZKHSmwfXT+uJZ1OVBd2+0myDmxYrIBTRwYxLp2EiJrrv31rF5T9oVRQ1m+NbpL9asT
euxzVKX4IvHbHKc4dCgakZiiY42kIHrEFRSQDeZugsX/LGjBmSi7pnxlXDFx4xxkfI7miBPe1q2g
OOp9rQGy6h7K69/quba/QQj7e+ACljKIER9e7cP8xr8CUEzoWv20mBwfSl4zK3/ZNlNpAzIptk8i
IFspw4E3eOO4zm5+lOYx7Y7lCGrGOOXaDshndGcVp7VIkx6QEenNPFXyGkQ1E7iglrijJN7EWZ8K
4+sKYWTCWm6DjMKtU6iZEzjPArpSwmYgJV207dIVAtzZ9+8HOwAydx+8NRUB3dktUnLHJ64HUOTk
2V1tR+PjD0dmO2o5MroIc2Z5Ebpb2+F7ohNAGB3eJPG8fzFSEXTL4yskFKApWACCdaxHTCwLR3vn
KJeOyvjrP2KzmZWnJqJU+A4rJHaCSh+ODer949shpIiYqBbu8Dd6O4OcEsqTq3vogikU4//DVBfA
G/6QoOk0EsRnlAieBYkm+ehX3D7Mqvwd82UAwyI8knnSDLmi4pMYOhQvuZ3K3WLXYeAkIIxYmypK
CjcVJV+vjX4TB4CPHSQ+k0eemDVEQrg/a5W+jsvBvGCn1zLdsDuWjsgdIbGqaJc+ZQX2Qgjr1SAS
+ASHLdctgJn99pNnFvrcXq8GqnCVm+VjhtN3DR6A0fzyCz1pM1WD+S5gCnMJPKUjsK5pQqLF2ZpU
K5a/ZA1It+BCu1vfYF1hpaSUhq/3QdLGKDLHmO8HUXnw2qGOihgfjLBIIFUy51DSsQBwdlHlkN4/
u6cgt+iisNKxztxMAfcBNMnWNXKPiYczNpRby7gg/gtLb8nYZuZwlazTo/Ndo2W3fMN9tgCYnXU8
7iggqX1Mb4jiuiL2qpFNzE4PQFSAkcsKer+KVJXcuUCa+9UiZQ3VpqmwflS5NoQwmU6vZSpUn4D5
msWpnL6gmxv4EM/OZHauRX3s+jQBkoSSxebDDjEXmJelw11b7j51zee4rgcpeQh48HiiJN3aVUNg
w6DVAel6CDRuj9aGhIr5yrPx8Y9OMng95qQaeEexZrZpKFesHJ7cv+S7rTN1w9QLnOQtJZZeZcyG
tFIMAawOvlNj3AjBh3Y3g4bpoFCg1znMlUzVQw1ZD6Zc1gxU7iZ0JKUcREooY9vFqy9mLL7zfInE
3Z0zPhM2L6R9WP2Ll/vlUl8UsMu6l0UEQLoMYKSlBt3gkcvJu3mNpCQ1hxoz3QCk9CJswzkv4ev1
k2T5ZyEKQbUGX8DpaMUCUDEoydeWGNLNDBxtF93UJYe2CpQTpeiTRE2Eni78utED6pThJQbb8753
ggLu7XG/cbY6KEZJwZ2DIBwhJscSftQJ/DafD2Tywv87cuLX48CxNzNSv8xiI1C8DpSgGAHANvJz
2LFryWPe1bDXiY0oPDAUmAI8ImUDey2nY/RXdIakGMXfGQxQlaS0Zm6WF5Y3CcVjS+Hp6KBSPcv9
Zb086j1vfsNhkSvFy49TocJe8mW5Dr5vcJqH6Z2FrU/y8jnPgKobckOHmOm5ktARwHXw3S+ELT5T
no0w0nZM446oVBPBzORwV7+IDUqq4Ai0Hictm0W4qCIhxXx3d4qz5yWkpbg/w4Jh9kgkjH+uOixE
wrELGSatDIr+m2/ASiUgOdKx4XrA/KuqSlwW468KHfBSE4VTaZK7hh2Pq+m9HrFhRXjnF6voc2Ba
d/J41b6tgImjVw0qL0zdtCk7EDT8MJqw7GLOwMNZKj8UvArZYb8AR582uIPjp9qWHFgIlp0pqOaD
xGK009eJFXoKdMNHHk7SwyCrb5x7+H+ZyQl3OurFDZYbjAJkpPEtTSfxOFVVgxnC0F5kfWZdphaP
IbeEFZomZmJ+SHJJN56fMwp/EYryEzvxlwru8O+glgXW4lU0cEQ7ZhQZaboZOYyF4V51pQkxoMSS
+hLvNhnxDQiy3NWIPX7aAOUUCE8EosQDZ9cs4R0OB+AoUPfKHQSip4OC0R4K+6wT8mqEAeYnKwWY
chOG2vacXr96gX0KPJS3R4WzGrKIXkWlvBk0oF5GykGUsXlQbIQxw5HP25cNEsewUZRurrZoIZ7M
f5U4PRocM5Vs1m21eEmATG09TwkYfjMJF7tpSKlh8JVHQ6HPfFvUm2YKOvy0tg9o/AseuuaLHPOe
wf3TnT5AOIMii9FiK2VdKXuWwUAXnDqDSgW+KkHlvMyFvFfKd9COB7rOfmRs9ODVQuLEk7wMHSxU
xBsGXnXrTLHJHHMD19rOiEKKwSvbOT6mWa+vkk8NMe+GXXbsYFNFvON/vEFGCEPTCBp0iMTTPhgk
WyaM6yltTVWB1jM1v8+4rFEVXHPg5p5kFbGDctK18kvIKkodaRFbj0SmrlBxdqUTP7k+nAS7jVmW
NmRy/kLrjdUanSYKX4kM85G+XQP1NgF5L8w1yn6Hf6RLe7bVHp5syQQiD3UttQguY5JJVvjSFW0r
ArLIyJH78FLPYayrTOIsqKeL6NZZMrPVrIao5CX4svO/MiyrJVyeQk1M3In9Ugt/yX/xErW0ekhg
+FjDeDEoIiF1aLc2wapF3YYbdnAKqQOcKFXg6QnsDm7xSUOO1Bz0F73tPqRA2bQIGxc31cjrAQ4Z
D1dsSnzoJhPbr7e9uzOTcdj5SU5sdyBJsYforP1bGUNzaQYL6it7aMLYUrTcyxNyoiw2uozcFULb
vsEKvXk51umI0XXJZBBcN/+0n4MYK5SGbXzhJ4ftX09JYHZjdcwrv1LIOaLB5zuz3TXZ93CJabX+
cHIXE0PDLY7MnQMNmQXkIpq98F9ifEs1hqAApJpg6lIzS21M4tKHCWxsmkL59oVo3nFWuYeODQL1
cdxShX2d0wOwaVpvl7urNUEi8PImc+7Sb3/PyEDfYUINGYXgPI76Uwvr5pSmLrRMPIzYzmZ4XJ6F
8ImAQ5vIh0nPhRPkHidR8hMEqJ9vsFc4qHj+WNLY+csmIRpdjXCj3zK/LSftwYewkBq8w6lOtzHq
Z9LrHIWtYFyPrWoN0ecto72I2DKvjbIry4fii0FubAciSQlzl6LPWodR23ZFFUhbvEOB/eeg2qLm
5eqSk7IZTrIkmI3koyOm9qRM4+ld6El5nsdJfuCILiS+f4giP18jYg6ZSwmp94KdnVhIGc4cbJSC
GOPx+6qscr3EaHxWpCrDZtty31/iBS/OYwrGD/IV/+z/w/vJxYC2ryd7VTAOwMx7ZDN1JFODZQLZ
gOxgBwyd1HjvNWLCaVu/FrAH8oMisLN5a2YF2OJ+C/BUjrYhUHboWbx3HvWwqO4T2/RAgnAvpUdQ
XttKnzRYSP4GvD42abEG83kXdlr3ZNP6gMiva6m91s3qPJsWlBS7M6qFAMEGKDX/RVHI8rKk0Sek
ZCgL5UHQA2cHDnVQWnaqWy+5ajAV8Z80TOtbqdVJsFPx8y8I5glO8cKWjEaDSWnW1Bju1nNT73LS
3Q6thLUrhmRr6rRPLukVP929slBAWQBDN7YLJvx2w5Cq1wM21zs6mBpbeXOHq4P4im/STnhp0XL3
2G93vGRBFgauvRiRZBoxLGXbXPLCD6j1+T9m/4abETeVgUB/9xPSl+8uKtDzqFsJu2kzaWP2/aWw
hODHLLn71dfOJEf2ZKdIxV3gGE6iHoUXqhwmvB+xZY1hPp7UQjBFC0mVD2xGo/j5P9xceU9092cQ
OxsIo75iGU61vfaypAe/lc4sxc+jl98nyDvDvSr5eAr5XmuKYlq1odYyY9lCuEQrEEu3wRbHnz5F
1T6hqdhJe7oL5/rw/U1CjlM+2ZFzIXNYXIUOrYIXMVYf1l0sCzDI9yL3Cp8ycqx64MSWBcjVXYMs
HQ0srwJ8JjOgEAzgPThrDw3Nv8b6dgBsZOFxpQ+QmpE8H46tEC/SP7KUvfoo3ZbaNEKKnF4lq4zc
XSRJ7Fv50PnJVnSd5M7AUtKS6eociB4JFFwqQpJh83/3sXo6cRAD1kt0zYvF0IU8eR1372/O1vo9
f1iHu8X/gbm1Iw/5ZfZGWHc4wOG4Ag260l4dYpkxNokAavuhdglEf29WVDSbLo2IYorNxl65X1Mr
uhZVe6ucI/6TpsBj82JlOfgNQtWl30GOB3Kuh30GPkz4yhUm0Tpd1gbYVNVocm/cjIZdVs9lJ4f8
9L8XEQM2CDaLPiy32rBUlHyEArRY2pJx/dY4McedkIX+Hr6en9Z3EODb0V77Etdnic8PvnaCj3BS
ELBm5scKOottGT2V4gW12bKa8wjcpI2TszXOGKkbBlWKshOsoIlrm924q9rKvxgjjDNOoeHoJeBl
FwcnPGa0UGBlRdPbdpOLMc6RtcSnMew0diGV4njNdV0W+LWJd8lx0Ji15FATMRL9I3I4qHyXmxxr
Sfmt4HbrRwMju8eMTBkxPMQsiCEQKweNMY8y9a/H0qeqzhmP/3d3Za8jP8jsBNwcOSUm0gm3QZck
Zk64fa0MuhIyq6nMaY+NXMyMHihnWPR4QCruH5QYmRTuKCgJmR/Lu1E6B8G8O6EmmphTKwomM7y0
ORauOZrEYjmfopriMurC58c0gV9ekq2nxwwL5/M/RlkJF+DZf4S8GLTQFbrHKNkCP1kStRhgA/ze
SfweMPNBOwoN8Zc2ycZRTm+cAbCLwfkrsDKm4udThdzXK5FWLx3wgzjbUoTzB8xLDkjHYBRXwkgY
48FlwWgN2RODR3pWzM/df/33pp7Ixt1L2humGhNkzbxOxqJ1JTJyK0/1MJtc364PSB4zhEpGTgvE
JgVB0odW2b6zZ2wrghxMumK106s2ReuuTcZ/3W/acdfbq1y2H6ZKUq+h8WeG3tEB6B0oB4brhbW+
SIZKhuuwAZITE+kdJKyXZBzWwAOYy7dNTqiwN1lQ7vqHvlWh/lUoVZAqmnR2o26rHgZICc97aQKs
gClb2DVpaUDNHhFXl6KUlzmgzI3GhRqNjO5TxK6CAP55E3GmK2UdpkTijYyrIlbMI+oZCEEFV6Wf
c5STOyedjR+cpJHQMAvjuH2E8QaClzp0FBXQBwdhspuBe3nW+CJuXP/QZNtF6Hc++U19KickOmKi
RTIrKDxD26DYKX6DV9ZfLYN31skmnKtxh7L71IySF7+FSccYsmZU8yvfAQDDSZoJYtPwm2Kdeicv
ClLFrk8xPVTdCb+564xPv3u8qdHyeIMkvVxllIIvGeTtAS+P9P7ah1uVNQfxWRTlWsLsS3v/mUM3
nw5lqeTvEbpwE/ioh+8OAgKOdJhfSPi+gJYFnHSkbHFKSpNx2zYYZ2Dk8WGA5GpuGLBObAGerP1P
pCayx76UES8FkAxrK4U9pb6f6MXmFY2MFpba0XduxJwIVRqokwHUBAaXYO7/+Au2Ol3tnfGxTSRT
V265n8H0sFnY26kQydgB9NN7f6RF0W+UGVtTmYd5oGBhSAUfy7QWuW6B9AiZ43eTfoZAyC4XJEZC
9Nih/r7cJl9OgRuPnzrCEGjsTtTw0+gyvdpKvMdBDA9JiXeMTGkXeMcf+OnwpVk6W5C/nwIsHF5B
EjECYkBuCJO1atCwvDIiTch5O9Nbsj8HYjv0dXQSv/LwyXd1wokdxrgsPIuWJhOJy2d/fYNcHN5u
adaK8gOlyaJksNurMWORWo2NOraqNXj0vdj3X7LUnGE3blLm6lzQ9m4+QyXx1KG/ya59WVc3xHeo
C7ENocomdaQX20f6/mAJgevGcmiPvqi73vvgmWEEim45rZT9wUYGlbE/hHkqoU0sA5pNpC+isGaj
AhjJiX3YOqkqZnXyb22KGE3QOlL/bHLEP87JDHDc0mRCQ3dRDXbOx2zMpqpAjot4MZryCcYFf3Im
wxWCWwfPPdku4+jjgs+tfJ2KH/z9cVdg74rnQkqNiGSzQvFr6GOCib6ANvGAuLV5zpRS29cO869t
HWg1aRMBolKyl00BoUg/3vKqSWH4LcnzsQQ1WyO2tndM2aUqXmcJbNHUrNqHl80egjv+OQeSMtt8
0GWyFPtritKT8LvbMYHKsbgjewrVDZW/Ab8HqhjhvU2lxkVmjrDhDfu1HUp354gUl7TEJp7t2UuC
TbohZVtOJtm7aCfbosmKIGcg/Cn3NbJKOvo8+LDX5xZmsoBJQiwjTqhFiRH6gJP0XwdWPRHNAPmm
zZ07YadVg7vjSkyY2BmP+JUcfuVFrBVarAaVqN3BSH4lF7yebA5D+VA2MqQGk3bdQqEUi1VRBv42
Ib3/xHN1LNjVN9ietTD1X0WdodkCbyNlizlUv1EoUQ+sVEha80WElXtpuztxt3S1MP/3OBEMSaFD
s51VlNg66r0SDU4dWZzWhp26eKsnMr9fr1r3yj/tp3wB8Q0cZYWIAb/GCFyyRKajqtq/p6wcLywI
ohIcVyiPGX1Jo7Kdfpw22x3/N+46A11tZktiMnm7cK8FzrARxNj4/U36UE0CTtI/Ht7Lq3U0Q4fi
yB0lT6KYIci1N3IXsXv1BIXIIOH1E0nkBXQ4p8OjZJ3snIHQu1GAD89Rw/70lObiix7guq0J6HYT
WwN/JWfLNNip8+hO2NzB/wIM4/uWSA7G5d6zFws6HbF8+LrcWKMJZRgxt6glpr4CF2u2JuAeGmk0
DVweBuvUCmOtM74hRE7Oocri1PlBsdTr6Er5oJP4bDznWFMmX61UL1Bim7nsh9n9Qqb1bfACfnuH
Isktm3VErQbg64TA2s8m6l1pPlvdfFN660Aw21+q9k62zEnNQhcnN94f6g2f030bPcnDMjlPOuSM
o8TYMjiNtVqK776k/r5cpzwd1kKuh6/ST/GF2wXHErWNHeKXCbVa0IjEpAt5PHgnVtClDIn2eQsm
TTWZud63E+WwmfO9EdRNkBLNb0HELtnYc1aMZGr2SFwm9ZJ8ayMwu0GczfDGPLKWgg7OYl7YszH7
WQhgwdTUnGu+m5IqyvmPoXXrA4gtJ7VJGqbVL3QIchs+l3e3RGA6p85l1OON1gNTTEgdlRfOwqnU
4fWAzdaG25/+K4shf9Txug/fYUS5fkQwmy8OKT0ly8BF9RA/qTXgUXfG7xMGcLG5EfSQ8ZB5a+1u
//o8EIYHSJKTCqTihF2TxEYD+3IO6mdOo+Zg5GQhChxs66aSeVchLtTe0znxILfi9nduljub5Cx5
KqnSDHwWRnzonsiVza0Vh/R4xXxPFyM6qakKebDGNje7QWjYnGfZrihVQX+N1oABniFetfqmIQMK
mIM7BAOLBTYUmPVCSy+LJMYxrbQiO604o61E/bSUaSTwkUtYfeBAyJLOiAnUoysWzEOth26t9Lnl
6NL+/PsleCLh5xQ6kaXX2xWIBe+xR+G7YkpNw3x/oMl+G0aHx/MM/KUemifJofc2O3h2kTyg+1ax
lLPgGr4tRqgxtl+i15WCjrp8x/82WUwBU1A38rsBwnw0qFUn50sRgs5Y8apojCrKy5j3apJr9tVh
nPpObMYDEi5BD+Idd9hvUe6XZb+OtrRBZj+8jIkFHl8hDJTSInmDTusbp89aUHuHsSyvumg7iBwD
D0A6i9WM8F7IyeNjJY9FKq+bHz1JufK3pm8sx6mmGxmD0FH+2dVC5YgbOVWqwKj90MJJk8ad/a6b
lpyIT4Cw/qNEcPUIsx5iaUvXbMvP7rMBSaxJU17ZegZLn2YvN5syH7PWVPA1a9e4HAfDQa2cmwA6
4U7ssCq5/ol03s1iGSuZRcTzkTW94BPcxwaDQ2PMm6W/D351MponxLOkOZf2s6SynNjRXESBtjsu
O5WCNckKvx/Etknww+vicR5GL9I9FkX/EHgfrZ4mv0fNYSTJWKiCykP9BNXqQeMXzF3UCsWK2OQL
frphmsVd3ectXisxxro0qjSSWogQHx+BQ5v9N62Tq9hyQPGef2VACKJ2ekj4e59qQ3f2jEAB0itI
Mp7qpCAB9zDfHjNLfCnb0m17W8dRDN/KU0qwGlXY4VJQdhp/MIfm3BRtFdYDXMrQqmiEsUMltBtz
qzKqEKicQeKJsb1H1neVSZ8AXNgKOHOoeg7/l5EprGXUjnHRONQPqUyG5sWrN0WBE50SypOUKRUC
CDh5qaGrJU9uJ09d4bYFRRgJs2CGOqyDPdsyB6gMfs7c3Ad5cfUcLOYtAYXDcHeBv3XcL8OM1OQQ
A3Cw4t2GVXhAUfFi9QlklZ5h6Zaa06kubCn+CA5GVkstofmlpsaUJD/qGBdeMB4Iv04UazPH+4la
l64kO7FqbA+R0EJEGvqda43Bc/6U1NTAsWVClZokFZqwYv4miYCZCFARj9+ELfz6BYAoHMjYUqMg
tIJjYjjDRUdFPt5S/ViT25m+kIAx4Kot0WT18w6E8Gw3xZhcdOZ6OyXaFyRxbn9HuNjx8M068bSf
p1FIhf7U3nWhvwyc7HQnrZKQX3TpfyVlLAVh8YXINqSJum3mIdBFYwj9AH3GQ1hLU2I0/pF0Wcfr
7M8T2lOskBgwv/ZSTa6ll9SlctG+g61vcVfXQfrPfjhlANrtNqXrbOoKuDaq7PErYbv3EjGybx8U
s44a0Z+cmZKXPoYa1MpHgUeb5Df7yaF015NU7v9Amc6x8Q9ULGw+74Aotzatyn4t6ocvLWYje0R7
V89y5fClgLZV3L0OcHa+jaM7w67RJslQhpkowMd1wlVmNoEag6JtHT67eN53lU+CFUAIG+1nXaxF
4QRC0A28LFKyc6gKQbKd0VpP8d0hUhVk5yGI2gtiAAv5lH0kzeD9j7gr/jYUmtO1MAvpbWI3OJfJ
xPYyL3Raw6umNjNAvybLENZdAzRM7XvySBNvFWBaOT7hc/dWrIO+uDQ2n6c6+EoHLRhe/vLsr7I6
x/cIZXwVcVKILqWAmcIVQp176OTbk5/ZJeQVzTq27Hf4Gh9E0srIxHhOKnNKTIQPamgCpg77pz27
O1giV2BWwYN6eOdxKtK6c6eGz0hJSj3fieex436ls9HfLch/MxVPEEUSq2V4lTJY8eOHibgns+x7
o9OBZnFXnHkobtEyOuO+rDYaQusX4K5Zsnbeb8wLIJ2XRgcR5jXzrugxfEODyuy7DvAJviEpUPiE
UDkitVWwKi+aAKKL2G5CuM6dC/uqoaBPKKmXSiMPV+uXaAQQMzBM6C8yLsPgEW+rN8Yp145pbbaM
vXI6/+Wjnfw+beQ7fXTZSjG0MqLwRWQe3aMiMY/M5/THLnzBSMbCjaox7SjtxJhP2YDOZGr14JLV
S+tislGsOxQuir77EggfvrT2rB7dpiMRmtsVojYLvmETWWnVpks3rwJq+VlkazAmzV7lJS/ZB9dl
hM66B3DtCfVLkWJJNMLk2hI00Z0OnQF56d484Pzp1C8qREVVFjuEGBOEbLRygmeOrSOAN+lLnH99
x7O1tKdieSfF6fmyjl4tU5XsGiRBhnTWaCwxgMdhf/2A4AhIxBjhXi/TC9NxUoRFx1S3DrImKDae
2xcc48XRL0Q+8j2I9IVye19JJ9xCzgKpuq4w7mxvYLGlDLbS+keYqkqC8rzXwQB7sxSkHDZWc3dq
UvhvlWkj5xMxLFBrsck0jesa99uk/wE8G78j7SgQe1PSooMFWeRKaqgwq2Mkue+GffygopbGyGaS
XFEdgxx+vnM+NyNPjjTTQ9CSyolBu53v2AHn/EXq1V4TZfodZHhcb2/nqVVXz6tz3LzhGmfbqnxf
vBJxhvWxe17L3hIku5Q5vh+pWYrPj0GP/SQwUSbQM4L+Bjv8X9TBJQXS/u0aAFBppDtvbcgziHXs
w1MtO7cHaFpZFN3yrAWOIkuWXIZmlqTcaJw8e5mUFLXcRkbKFhwvGjYvhL7GECJMQaNJ8c80wz64
sMWP4h16klbQIPy2JLkcdNLT13xj+b7dDCLfDKkTluZ4/9ooqTDZ9ZXyl6nZlmORlVU4QKW8rdDX
zBFe9KACZArMa2TCXSd+1MK1WykspNkjh+9r9W6eFtYuc/m3e/hRO2UZ0O/7mx+TcICXpjsTS6c7
XkKUNj8akLpuRZcsVpylIqXAuxWkCNqVs53iFUq2ce/E0De7NSOJh0+DPcPPZYgIKCuTvf+8lOtq
6Ksk6XTVErtZBaWWYCz9Sb8vy0wg4CGUVAOcBTYZCzvIMolXgHXXT79Z4F55uihwAw2hFKtiYGK4
yaE+LqL5AORmE0w19+69oLweQGPOGMysqozbi+0zcy/NJRF0bOJiHkVFVf5cVkLsUxF5tGtdZAlp
cC6kuk/4XNIcAVT2/qr1jz4CQH4goCJJGdOco4U8ToL17vMkw4BgTWPuF5XIBkB00lMlhRpo6U/H
G71iHChFoBotjXz6aIG6nS21E7vD7HfdAxJp+/Mu2YCoLXzKGyOCPmrwWrD36j5fYLFdncoxb1yb
pz43/OiLnh8s88QHJJG7d0mpbEA2YVmhjJUoPy8cL56eOqHckQrprgMDR1US0lH4nHF7VTYtu9Om
dURwrTuk49vgrqnA6vv6fqmAAjhJp7K456OGgphJWSoFKIFbNsgVb2KSP6gZ1GC4Q01NSdOK23rT
Ty/1cqRgWZTVrSmeUZXAjhdD0eW/NFvg737BJoySMGi7pya8JKgKGKRFncM9X1J5lGkO7kPsOyPT
2P8bqNmeakhbf7Y7LZe/WWPkoWHIivK8JnHa5F1HcxZz96Q7szzOM5qRh26MlR2Wys9XclhWnLPn
MLzEjqcFykL+OeMSCwdPs510DBvr/HkgB+BanB49msxbI1VWfrnho6Vf9eJrFq2FuDdOXUtgN1A7
HA5DC/Ki+ttLFxS1dLWIxKpwk5E8CUjh4vYOVj6Ztwr5wISaMfRaTSCZf3g4uAMSmEqddFF3SEGo
B91cVftgHW80hzB+VFJ7YkPXUSs9B54zq5lj6evbXpqtWZknh81IC9pYkrTEXOwMMIpMz4q/k58n
ut4E0vHdLePFhQO0EW5qNgiEjQZmIJUbJzqe9iEGq7ym3ITwaMTOz6shCsGDSUL9y9U4vpTRVsye
4hVJAlVEFkucaWunI7SRlOldQyDr4RzjHyvOv3sQB8Ok7zkEXyRjUaprOf2AYeopxCQyjsLaexQ6
3ZYRLdmoD7IFiFEGkM9B4HEbYmzqKXGbA6f0KZe11Pjkiu2l5eLg55FWWARhj/z0jUMovFolmXBE
OuyKkD8JMj3wJnRBwiwEtKMzbnilZhewlNqsiDF3kV3YgAxwoW7ZNtEHfFuzLtfaZY856cLNJ8P1
HJTqDpa9h80C4URd0H52Z9pmgNOUCkYZNYQLvr3ng6SsdaIKlCo0PlhTwRvKfFooH1qxZCcThBij
bfBRXmNVPJHpUcCty6nOIEx5bFV/rI/mZulZLgWcUmw9xtXF+6aQrO1a303Ixwfgo6wJbgPny7ur
yNVhQRB+89HiHjH4zrL96pZjD29/PWMl0ydVFxkRa8AWD7lg06hEMU5ZLpsXEdVT54xnmKBhLxcT
QhjAq65QdZ6XmpskHOkvedT6FasxJk06UwTIwdlZhKZ5Zh+auqTgXUlkYs9mfZFfxldMeIwZFbrM
604s8ahyCC4q5D21I1dY1XAkTC4U/shW4AMKHvvhUAqwPUuVTCsjdDbHv0okk9gYE2YIsQX/jQl2
Z6VIGAqNysCwtHK7GWmlVGNkraVGX/ictI1L0TSKDHonEsW0iHaAoTG3xyzfscOlx+H1wyOTKpai
1+cJ7LbyotnQ4+s3whoL3K2bh+TB9qolwSgrXZMaDHTH48B1GWDYwwSTVmN2X+ofTf1PWtCy1SaC
/497kYlsbaqy+CWMtZLMmVoH6UHMrtPwV/nGsd8bW/TwosrKTVQOlXfP0bZoPMEybVkhOHCF45sY
H0wMYc+5bitmeNL5MwfZn9WEMFcm1pnXlXVBSLMuX6ZLO4BbHwBpcXKynNa6YaaWfMVYeiBZ9z4s
pTjJt3sM+jKw0iSIYvLn91KPAXexJ1cikwwlMw9KDUlAc3uwCIr/z39fG6cIj7v+//tz67Zx3kS7
FrefEjQIjKGH41H2M61xj3rfvlIwKCkZkNirFOU+xAuEiQg73dunUKPIOKwNnLhNGi4voRdLtGL3
zBmH05BMRQj+pZ2cVnZlL1o3xSzA9hV75ykPVYx4LWGDNJJVFsCnbiNsMRn9GKaLbE/zWywQuIBP
N4FZenTB+60jR3yrtVdXL2YaMgxWG+2lr+MuzfhoAXSvBhpnRt2x20TRcBLynIzHK9nwLsifnBwb
VL9m20ah6u11M0hdsel6FtYFtrvlNef9AWQNjWtmJbbQV7aViR8vyga4gha6/LnIHUHsIN6wsHVD
4jk6OuH0lZyKVvejf7LP3rt1g6ZZnkV0JQU41VwjVd4l1FfoKrs7lflvPQUOkIvHj1BQKWRlSQEH
VA+X10WS6WHp+leQoar2ah9LHWtKs3zK15hUeqtUsaeRoUKn9/7gaLXJThzEfj/H7mDmRlNueNE8
fmZL8ojXzfut5zNJjTMtKLc+aW60qo+1EvQtlags+WHAycDhXovguRklBcguJpgoZs5zk5QHJfpt
ozFwdT7I9s+0dlqW6WK7EsGZ2mNFA8JzbzqQgW80/lzs4gRVIqE2Bh6zqgxvQFF8lPe06aQJ3KSt
uC0xPJeCyCHedr3XPKPDm2GKmmseDs+XIexk4OWOGF6HqeJMuzYyno95voqkYZEKUi2uY4ovNRlt
ZgquPjArANs5Lx8KM4z3RI5MoszP5M81I1AzayBlEpBRY4ZOEqVVD57X/ZF8lz0W0eaEE6v/cNU0
7uX11J0VXjDFqLVwlu7bePVeB2Q8YZunAREjnj4imIi0r9kbLSrTxiuazgfpv6wlJQfRV5ab2kYl
DGkltlECiHeD+V4/X2eINJdIv22geCqtYG/DKxwRj+/HYYoFOpPWANqtwaqAwixczGkgylJQZHpX
Ij9zGkIZ8sehM2a86iggQ7RxcCDjLPAZByA6DReIK7YJg87eXONEB5JO9lrk7nK+W50NYW726CGM
sQIsARksrU+MCK26nTsnX0M+ioiaVkyDom3Gq9UpH0HkZJ47VwE7KNo6gGPEy5OTCP5LYRVUmdIs
k8eOcoPnEmEiND7Sys8onf/1HKuIjCqglnNx8w97MEnPb4xRgWY4uGxNUYgVX79owy9A4FbrRlpc
Ng5IMq4xOggi3kEOQYYF/jPFY9NkrNHOjauBuOLIlgbc14dGZ5mpdwO6hIKXaO7CKoYkVjQOlonY
ryv2H36R++El0znt4gHmDJ881fR7rKnONf3qzRe/Zl+gW+b7eBn8oySO9diKuaOlROPLVSbjXk8S
WAlk/tsWMXqRMMH/ZqGPWL+YY34FiPiVuvmy9e9zklqoXOyX4HLbuh5KQVKl1kj0j8GRy789GNtQ
sNQELurkjfgcCcYv/LmSoENP5dw2SyNzHHIR6ih7/GGEE7z/3tqgqtSLNxIj4hfQsUzG8fkrVd6J
TPSiL8ztv6U701iD+FG1H6IH9tOFE2Jlsjc2V6H3mRrdulkoUgLuC6iwDLBU7Cv7LhQsD9qsM4u4
A8X3wvDT5l42oYQfTpBLa5HN/54sgB8vhFtEvVtlpd6TgReNFlcN6QXrH63306At8z44zb41BdH8
nc1cJB9M43oksxQgUamiSp+9hyBPGrV0BrOWTocjWnfc/dDP3vdcIq03w7jyMfsWpa0FVvnwLQtC
0f4xCkUNagDTfw8NfPP0BXha/Mips36R6m7Xp7tWihP0nX2epP0zezwBHSqVx9fauGBp7TWSDodk
lIHiVVmUXef5F+wlg1Mlrd4ArJNUK9ck8CZzgnlpw5hP7/5B0L9F+0S+0xyr5637GlRnI4rziyV/
uL0MQVlKZ1UXvYnwI7ZNP9E3H/v5rDPEzd9+hEuBq2ofxA7vFanfTWtkyajBFf8K+O0chrK7Vvbu
KLNnJFfXnnJAWWyKoaxo+O/MmuoeD9JKU4XDSPMlHqN3hfgKvpbGLgh6QTCFbX5xeBrmbjUhmD2H
JyBCefu5tQiPJsrhaHiMjJ6JCePJA2paETmxRFtFEEF8pwiv+zo1kjr7wOmSeMzShfvqQZc1vgG6
Hlz2ZQ2Nb4FeMqW+YwLjZDVHLJv7ij+ljEnDXQjJ/+fjdB6rsLMGED2HTRQ4W0FVIPHgGzaHSDBk
1TeRrB70HO/5KmQjWPosdj2dHW2rSASnebyg74YKHL9GAZq/SPjCGhWcVpG0XseX5xdT05rhZG5Y
/dGCND822vZbyT4jTuH54Gh1HGYFnz/t1GaJCOuhaWD+hGnUTLUGfVLZmyDx/qYHIlFaUJ8ugrIW
ciC6UWtY+NvfkUGZ392e9xJ9Q4JhNot38ChAOoi6aXbrY/n5zpvdPgoEi3kD4ilI3W/G+Gn7NlKZ
BnMQQvrRmGKA31KxY7ABEn99QlbUFPvqHXotAPUPS4Ha+/fKqLwEZ23cb2K3V5ISDpZUL2g7drWE
fVixXwG8/HBke/nwEw/xNnBK5Y0nQInf2vqetZNI5eZ+Ib4OIAKW2IZh6Q7gfQcMoUoJ4/S0hzBJ
yG7NTzG22OG1WOAgQzlNOD41I7R+e1J+7DRIl1YKv0FEXFQDA59xZ1E16S5IUkppoZv6QIx5/TxX
TzFMj191it4KtPyJhmayvgF/1I+a71uQhPeJYC5XftweM4pxTgXPBNTcJ6WLc5mW03SHDeL4dtY0
eqzQQHIDtu4/wdDqMtSGTyehtfH3aFmSZGhlq1E9GDAiG8GS+hI5Tuo6Sm4fvFDfmmFHTL3dnK3d
sdApmZjrlE1Na19hFH/xSTrInCWP9MSHBBTm46Gr8MCjt/GaLad+N2SYhUEa6CtIvmALSECboJrM
QED+Ao1EVblRbxnEB8wCB/m2cGZOxuSKZ32Xq5mTyFY8Txn3T0OxnAOJRr7Cn9hJHkfTeYUevQZg
hBCjDKLgfUnnjrI+FXY+VO9rcgZlKNu7SaMT4BZi0TDahbwicEqTGh54ry/TIzg9zx3Xe5l/HoTX
oZXZ9eb3dckqWjRYG2SNvad2O+3P1QYl18DcgQGvTpF83WpyO8lsJIVVeXNMPaRPhtfgCPfY1nVc
c+iUMWeLZKtWXoODvgpnc8Ay3k9FL+TaWq4TksdCP2qe9y5NNHJ6eN5ia5zU1FWmzY4A4fZgiKjH
63viVb0Syk8onHXeHCp1pjpQcjmvoOmfYFBZdODI8aOZEaGCneUJQPwy51/sSF1Vf9gCe60Bwkez
4xLPNDnV64WdKN0iAZTPWQCLBk2dE34ZKnQg1vuYHVotbRCSUHd5Bb9AJYyTQL3Z1n5M3khlce+L
7WKvhwjqUbUAAqScw4R9zSeiTP/QBgImHmpgjKc+LhUT9X33vIOVT9cOpRQCiz0BXlLwyrKJfJtq
ZtseJ8mXE8t89nlCl0PnDwCh2khf8QcylKeWPwSwLeL/e958DHt4jyjtuHNIplPoQkepxCXJN+NS
IQGkypIaEURzETMm/ssaVrHvfl4OpaGndJIYnlTqMwu3K+y3dUcswcz8FAm1Fm5bGCfMN3BV3HFK
4F6XlXjfOGja22wW4bBdgiTlqa1upLWLemU/+gJ5xw/O3jbjXOESHyUmd9ro298OH8Lhz9sFhLPa
yoQLpKz1cjIEpDXX3+ncTMYL0eMzUSxLQv59v+ybrQJIvUQ4VKYJcwY/mOCemd+KeHfU3Iz+Om1C
VWlYm9PJNyxkS0v90WUXLrM5k9ZjSdm2KRVo0jiNGariEiTgUYiLMbnN3yy57Ew2SD6wV9RwmSog
6G+thoQGru6ceRUmB3+KZYHv6LgrEdtpO+CqEeEXPZOpxfJhgMGNtPEF3v4XygSRPdYse1AazOPn
drYO7rx8yHPluLzeDvSkL3S5FppU3rRQiWDJKzUp+3JSalhiXzrHTbxTcgni9r4cfO9lHCfMyt9E
UNW5PVz3UTEdnyFQuqAX8wuTumQie5CdOOai0qRjBpb4DAKozhd75ptA8yWvBwavNA1XTAu6NkTg
Pnn1DY8hAy6FRKWXEaO4v6ice5tSMzdFf5VGqKnc4LhFbv36jz7abS20Dbl4rbE2FvtcXqPFwOy+
FaM5gl24lfzZZJ4YfkqFZMSeCuk+6UECVFKI8qctPFLLpC52CrRWPSZ5pxSuX/RZ/i7peRIZ8hob
Buif2BT/br5a0f9nkhi/2YtM0lZebDurBiF19kyEbgWCosmDXk3Vm3K+Kx0OHWC80YHwAxwjCS+9
9jVwzRf71Q5LtFBk9JMOCC0AyC5dFEM0ivd/eHp8btBhdfZIN4IpmesnlaZIm+FbO/jtYUfogitN
8Z64cj8Xl5OUG8XWq0RWWMtoLt1wD0XV1mC4h8s/DABHvsGEJ2mWrkogbB4sIGrKwRa5DnX9ONUS
ZTtKY42tuPLWY6qmtDIiHNnhTxdfRnZLCB8mdjkT6ESrHPrWIHwmNKYBk50QhHW6feXr5aBAXClf
uzeXDtSTFL3tIgT0ZzMee1KJE0OIMQkNlyIZnd3Z9yxkyJqLbN8bsCqUWdyXXgoStWaKDTy8U3Y3
fESCr1Llo/8LnB9WeWr2tg9IO50hDTT0QUyDSBTjl9pQ/xb+VY/LaFj21o8puRNblPSOcIH8/yAG
ovlr2WrZnPYeQGFsqtZgzySr7bn4SLFVLBlv6OKnX788l4UxSahiCmDLJs1MgGbWkNL0pzKMhBQg
HoLvZH6RHBEun59gmzP8eq+VsyN3rNVF9Hg4q1MbzZMzsdcDnNLiv0SN3auJ7aVn16DQET7v4oJ1
s6Ue77pp6vpWiHxMQL3bfQUQ6CLxSMhC0znobfUhfQS7oXCaKOWs67qs1zkoHs6xRi51yWzFZJfF
ymu2Lz9oU6xLiIMXLhVyL1l7UPQgBpcOYhhifQP9RiitIrrGXbD18cHiB9CwqujKScIto5iTRqIe
ihXVU8hCpWlZHNR5euh7AFm7l4reYiSQdpWJIm6igWjrhCczp0qzpkYe2O+PoHTL9L0wvh3cVopx
vhPpe/dxINZWg6AQZKAsTQUJlNZvfaF9v/INtGAq5tEk323fNiIfSTTIe+A1SVRTkx777nm7Ti0d
ZY5pie3I6d4fYARVr3Ip3pg4IkUsft2TMk/QLrxQl+LibtFif+1pn0HjsZ0oYTrP5LKLdrmG+qyl
CnlHdsuYLUF6OQbR4aXvBbpJc219yyRFas35lqVNVDWMCe5EUaNhjAzFkzI/QOUW64f33B5Ec8Ch
pxG4RiRFKZc4OY80v71JlEaoK5D4JW1eOUxiYHHjGH1fH+EktIox17kIOAnpDS/8rmRSi72rVPeW
wHss4vB8HGb6a8+Ix2DxAsKyKZc+rnY0uvLBlGf+JNOK17ISG6IAmS4OJsmVUDA+K298xkRDy1ws
z2V2PcXw6ZpzGJTPOWQPFcPrc9nPWUT/ksnCSJGzLQhVwnYYBd+s9+NQ3mSKaaRWzlpiHEfyeO/m
vzi00oPon6RrcFLL4UQB6Pa/e6s7J6YONHwXxWIvrEdpj4S59hpZWABqvZrVP6X+swUo9vst+qB3
5I9kZHCDmPFLQ77HkivLThRD5VcQC6RBcg0Pl51wXRvwOGYW6Arcb5adZ1UDfisSVmctFwUbdDOH
UAM58r/VhEhSuIUUVm93masQW9LBmt0CbcP/BsAZ6vSetbWuMe7fOXz3U+AvmDilm2pEyQZ3Yngy
FQaeUIm9rS6EMvaEWtGvvH8uWsjWlUp1M+9kOCPPatCxvjitzcOUPLfh7bn9oHKItgKy9Ihx5qas
P7qZjX10sQWssTTsmdEszu04xVXKOStUvQwL8Ix0gFfMx3aCdy3MkStqiPpMgZjZ+gSbpp43Hv3f
Zqs07iZsRJjTW49Wn2IKbUM4AsySYzKuvmoskSkbioiippEVN5N5kzR+P3w2PZxTOiZU4pMPCey8
/PrWUvkwNkUxd7FpMj/I3DjNG8jnVRfFXVcaZ5V15fuLF6AFso/2Fjxu6sAiblG6k/xcXZype7M9
sa47RtsrRpK5XmA+QKPRvzrC5RY1ROlT5OWlp0KdUYkfmvp5t80i/VoWN1kj2oG+H0Rs39BM4LX8
ygmaPU3s3oevhmG1nFSA/tjYqkmETL0bluOwXG4b5f8JeNV9BGz7C0hfMso3BA+WjFVZC+V8d8PN
rjYzq8COrSQFueoXRXVTSdPLyMoMHL61treq9OVsZOJInBniCdZUHO4ZIicNi9ug0mTZ/V4voKXN
Todjzubgy31VGOZp1c2UZemGM8DgwxQgmwTEnPtWLCIsK7yjt6wnwTxhFU3gkW+AccDMXcnegn/H
IEA/EVNrNlsSt01iWQD+HlrcN+aU3bE4U1c8lZ3LTyK0+K1DaRB2bqaQ9RFH4hGWHIUKtw6NqWe5
QVUcby7rHjUff6DE6Z0ZZv/0N0KIBsJ/0lxTlCRkSuNmv4j2MOYdhyhlLoZWFiGvshbOI9RXFikW
o3WbC1H/Ult58fHX7aQE8bqjQMQ0AJQEnSFg9BYS04MjJiGuvUX5w9p8dtnKcd1uHPWo2HoaWUEG
dDPWCdtcN6GwqLkC7T/44FlGP1ymhbDjOolJIfFiD7qJCoIvAIvm+doHjZTPw5jtP7GqZsg8GRZe
XE/wHMGZO41RpOQ7kDNKYC1sQ+/8Cjq9Js9zFU6wbn3zKC7f5dDk/NdjZkjhJnsjA3L3Ff7GJCX6
evJkP0uXTka6FgtDo9jx53oWAR/GYZ0zjb0mEe7rWkxBV/Fa1cKN2WT6zlimHfVzYsHz0iRZFoAB
F6yNEcd/acpdKjXhaw4cU9Tk2IdTXeoZToAHu1O4uNb+lPam7nRWW3vRQ1j3N2Uxj03EFMlWyjg3
UlOWv1DaDbSTn5f6wVU5RfIHNfhYzuBqYu7jIVByGv/EmbgpVMoI9p/lEkMdMI4ZtJX12Wj2xhq+
bhoyzLQTsF/jEitPd0yFlpAQMjMs9dr8LOOtqLk7IYTm4Elqs0uJGd4+qmq/c88Y4vqLz5PHXyev
kb71+6nnvMnDUktM3TmzePa1ylNUTsgSUDgmbOKIZWNrezGvqLzSsz83jynNhb55csrZrEbjWPf5
OrGriSb+gpStN+1l5xcSzmA9JmMdpijdTlUv4OMMmKQ9bYtkiDqfWaJBri5wERWeXQFlBRqmo6Ue
VMFONZMQyDKFARB0Cfzdz3wAfzS8kiAkdZJIub8+DJiGczx84s+UqpJMhpgCrU9O1FxDbl7uDp1T
vOHB/XyLz48O8S8hfNAFaBqvGRoC/i3pnGH2ofU0YNJy1bP17yIHvEg9ABMb5RUNUQNeEgo6L83+
dpvEao6YfGYsG+FRP2No/97TDlyn7VmasbmOttuKR/EOHeydeto1mWoQYSjLFdS8uGMfXxPr0x/D
7YdSug5pZVGlCLhgGGieQnORLgHcwTOMU1chpy201xcocpTZ8LImSjrO5UXkJzjKAHU/qnNcpL9T
KaXiQumYf9Pd5PtiOTIRORmNcMp8Xqc3b20o8ZWyOp/UfXfG6G7Qcl2EuZOqn1p7QT4xWDe0Pa34
rWolBhebbJ8u0TdAxUTksfYMLzEKDM7LicueSl6/N9ULKI1Lmi41j36dk5edTkfpS+RtBBSCu/1n
qZfYd4wlx74OjOT256u6yJpCCCCb5gIMUPhj9e8RKxgqjlXZUvTnasMb9dq3frxvcFu6R9WmCZrW
Hb4vH43L3P8J+57r9hOG6FJTFQwXM5TrqlC4WiT5KJhmP735jd3QnUt9zxqS/nwjwX/7L6WaRRoi
jDCOXkJw342X6q6a1QFHznZNmyCzay1aF2xdD65OQdtqNn6QW5LQpA+CHxB4gdi4SIKefPreaaOS
IR9bQTaGA/12zkpZs76FHlzyEONh5uSa6THHQ9OYvjLZ1Yobpa71MS9rC9rtKefaNfei+mRSca/Y
p5YBc8Sl/aCoKXRj87SJim/BDVJxk9LH0xbxIHJvIqDmJH8BsiXCgzaE2FsJEiKLBCfaZexCuk7K
4v/DuyYe5nwsdZ1c7XTeChEdztcnDiUOgFm0aLbx7OChIJaxnvmzGprxRL97F0XR23DGk62+G02H
kSoSy+DIvx2BxXOzOvNIJiq6zJ1oiXksqcjPCwQo47hEK+PqqT9O4ycdU/xdhvZoVYedEQkFxvty
XAycMI0qZOdWaV2T3AC8+vwjxC4+ymFyF4+KskqAPKOpQNsFVZQtlMigRLjDjxO2AAYSNDaanPuJ
bYACt7MHOg206PmnojipcbDG+ws33xvbVfTTaVssRtAVhWNFzKJQPXKcGOk3HCLBs4Ywt5fgH8lN
MjYGlmlXmShjV9Fr2Vtb/hCAKEI1OR4HrrbkYjHD0wEabjT/oV5oqFJSvlRBNbhpnZ/vQBJ6YsGI
LnyHkw7jfMOQHWPwpP0CKMO4KkjbOBdW0/0yqfEuQOss+GkMvYakcINySs+fz7hdwcN6rL1mG712
6sJV7W1G8Pyfm0tqubLTnTIt8tFfzADSSUBQFkyD9/MufD0PKiseJGtusgPpqnXVh8Hx5JAYBBXW
JCotk78QGtDSbP5Uq85+p2zpsW7cM6mEoAD4MAIMh2jW4IFKUeBJHFhlwLWJtfhZgnXCKF/bnsKt
6qa6gJx1gPmAW2sKTboebGUnYdn5EHO0/WsFbUAlR2E92yw9rIvK96MmxCEQj3gqc9TsAl6Uxxnl
n0H3auwdN2W5ULV53ZqsYaLG7S+inFl+Em0iz2Vjq6TBm1guwISe/v5/keoiLF113MRBgLLYKMbe
3nqcXCsgxSlGktjO25FWOQJ3FjFiRPb0Iy28/tTv1s9diS4s979W5Cc8Z7xd8j8L+CC6SqVUgUON
vVhZG4l5f3uqwKWh9F4oxa38NpU+JMwZW2u39wMAot1IgP8r0qaTMcVkLIYcafoRAviRoYh2YWM9
h1Bakke4saDS9WS1Xx3IbtgKueTrx/Z3BhHYGBkj1hBml99o4PMCjyA6JCoE6bc8HNljJU14KQYi
cMYjtPtygzb7nTisF++tL+30H+UQgndBjNrxJ2qGGAuJx1ulcHprnkbuC56dfZC7dqVy5oCfHe7g
pvfwmSFaRbFpoK2ZYA4NE5glrecwazXn8ejM0Navg2xRWgcBMRpd2h9hF3aN3MEDUBbOR3UGt4cQ
zxmj/DfOfC17m9/ZuqhGyxZKp+QnPMMx8Q9azjFNvds6cIr+HUw/+dW0DNJ9bCCV0H/o1BQgI6YR
upHyMSDBjrw3PKK0aMRdVxp79gbOG6tCf1HADKuLFKMAE2o5kYwfUiDHSmoAyn48RcUEmpbGOuMC
QLgOUpiWfwROHypPWbgBf2U0Mw73bpGhYYQgcJ8Yczh9kw0dqu5ajPcP75kPGN/BHE6XKyA3NYiL
i1qYmVClehMVDF9Obp2Sw7GSQDBZ10Jm4w0Sq+MPfyLyG0Ek50kNURRsqc0iqzRQ/z29tm1z6AFK
5oW/v9CZqK90a1+bNB/KUHWyak0iwSbY4TS5bqFV4KeOpgmjFg1x2xoDmu4HffYMXsaL83AU7Lay
rppJWFg8ha6gnhUkc5WaX6JUeWAuZHAiLO5rFOtuUWpBYx6FMkrHA3zUwfwIGtWlzDEmVurq3kI2
jIe21r7UlvBZHkEN+izIgsToFgxNczIRofPKjTlWU9CTS2jHw1mXoua2AYCkQorsO6Ha493QXYJl
bsO/2bYDd+zHZSTJow/g0Fvzd3yIRUSzYZCYHuz1LV8HN4tWqys+ASY1ELg0WfdOiyLd57eJYgTd
WZXFpsSRSY9lcoA6PVukpkMLm8pr5iKNB84NzT/mEpYgpqPLW4BMQyp9bi6bUhuHtoeQW1cHNERk
zsB+TmW4YMv086Lnuh/gK1u90wdGGmRz86+inDhiaokRyXLhG43rxc10mOoMpC2EBf5FOkWii/0N
mSeyxeW1q2uyicVII1ibN5TwWyQtejzITj98ELvfbekqglgJLU/eE8yF06hqZvO06HZYTmLyR/2F
R+5hXoitr3kslPDOUHmTAjbIyoxOB9/5Mg0PtiwsPkY4dKryja4+nwpsf3ahLxVtkhaA0yKNOE62
1Zg5veRDIa1D96p45YY0khHknc4h/iiHdr0PRiEnUzg6pJLJt4DCmcRE09399rNNcejXdIGab0UR
P6gPupKXi0c7LbvDhrC7QyLO1Qh9udPc8xd8ZwMd+/CviXpOOkO5GSu2kLmfHHzVCqZvYdw8GieN
4LB6yxvLaN9FEHVh3/nMVYOYRDsSm3+TA5U6mnUjT4+IigOBbhHOmyB9kgI1UDBK6iKKEU4/8ZfT
/bUT76xhEU3bHu/di3WlGXTR1xB09/QJIU+TC62ATz0nvEC0so5QxEURQQIZ905qqHKYIcS7YtdU
QHFHO9FyM9ARfEqgPG/sMpsnhGALKOnyoFGU6NPhLx9/Iz9Gs/ZvBJV/AnWxpRfsCpw/EOqNTRbB
zC6ytcFhHFDizTs5kF2uMqYKK4nXH6eCOTaBAZFbn7x0hkyMSyMR9H0zaV1+yaJrdSVnqS8vc6qE
j+75isgWJMtSNxBTm+Jy8yBgXiH8CZzEBlYJyHBU8ATmwCqIiqYea9CbPrNh3EH7H73gv7Vuy09j
P18hFLYw4IQphTGOHyUZxuwGsejgMzsH9cwALBuuEMmNfWF5evCzIjQkp+8GWB/5CmqucL8FohNR
KXViLQZGh1uiJq2NKnAve6ErypazYeDpUi4cydqWHmZKmQtucdNrfa7AUjtO0XFBCDXjdM/LPv3H
ya927qy92Sw9I4K6DGJvr53lfsDp33L5hrSNvo9cDLfB/L2OZWrOl+SWTLwOG/FXZYEopF9gkS0z
IT7W3v6b4QMbw2mS7ZJFoQUshUAi6SiLofP5/oTlBpSEAbZwlTg1q5Ji9XJL7QBKQL5Alghb8u9z
e5hOHK6njKrlduYkjy3YingM/xm7RKKhJZ+7uhBb7lPJuVNcxwCAFZfvx7HSbvsFMX5QOHU3aTIA
tLvaM0jcW3NUq5Uwb+MBFL0f3jHZQUgNoXD/7lc9zq+dD/slkhiszLXZtlpqqkzZcDbQrhxNttRY
PIMx+9HPwapogIFLJ/NIsOhikdvCKHn3UpZ20XDvxJ+hlPryyCzffJXWkeGgBaLNOKixoe3tj/Fa
ouANz+/SZcok4yA29eUV0XUUl1F/UJ4PfhprdaxPEA5iYWnYI5Sk29WR+bzuOJr7khQ+dG0jqvci
UQ8yU+KDUNyBGQXai7LCXPV/BE5f2CAtuj8fkGI9KA5uq5c4s1MTb64IIt2o5LSowo59W/8zg+R1
X7h0e/t5XctPqINX2E+7w9hhUINK85O6kxXfR8Fn+ez1xXbIUlPmvfLyQOCLDxXOJDD7+5d04NzR
/XxyTMvhre+u+3RIMKFTI+NxbLNwqgBYnVsgwQEiwA5FNqoi+aucSlnSdpu0yFzwaq04v6pmnnOr
mISMCiGxxO4N9VAGWwLGnXTZLa72vsJqolFzx6BiQ2NQxbuVg6BzijQOvbtM6l11OL/G6NtLEhUB
j4KQwZ+6P6s+KlDosyucYGGQqiUIx3pbOUlUzfw+uLUOrko9CATZKOnkjn4AP2+DZGEWd+zWQmuY
D2zRf1jX9KdeFJHi19N2nM0XZrh1vCr+JtxhkrSZLSti7j2RiGQdgHkavgRyfwJkyIDAx3+iOMzx
wvhIZF7giZKPpMngT9xokLPebtxXZAsjgDu++WJGy5JFuKAdmNOoJkwKTNbxwNxkkle7hQozHAQD
WGU1cxDEjBRHeblA2cGGdeY903J34dyqHvDREKWq9QsGB3h0vAZWVLkwMEApRaVMCJqKxzCx1h3I
BF3RfieUxHEexuXFyNRNRymYpvcq7WORFJ2W961kcj4y5dhgDSJBLpNkMrRC8O2GHkxjOOCUujue
7cyjOQTqhP2FNJ2D+iCLyI8LyHqAbHR/kN/LcIPGCKEYLoqFA8n+dpz/+O3vHHDaADi11KyBykxt
uLcLJ5r8RqWobLTFxnY24+s/sknBiUSVtHkY0Uz2C5VSFLc/0pGpdym9yi9WvnPqnzDkAQdwjn3r
1JQ6JfXH4arIp8R+77KMNTqsnO6PvogOGc2D1UjxooH9D5oyfuet7b2oG2tt1EaHN2f82mibbkY5
fzj7lzBNZZhMe37MfZi/ITE6H9h+7O3n6d4ctlXfVAlKJo2GRLh6k8VQAg05v+L3zw5Cw2VBf6nZ
fifD3Svlzcrq983EN7tr2yH5BI9Hr2xDKVuR9Lzl83V1mhZP1Gwl975gLMJxpae+MOdo4+uyde5T
22K4GD5kX1+cW1sMAv9pG09gj9BTYrKtTe++c17BTcQE4u6taE8sCfLK7y0586zKgPZp8lWbj7M8
F+AA2U37vOd7Y5DC0gpqE5bovnNF4bwekRi0jVWGCUe6X0LBhNM88woG7GSKp/WWdQQIh6dG+sgF
F09qkNiv5AqOISFfg66racvbOSbW7avK+iN/Cvbvp3Y6mrtbqqnJRpcyru4A8KMORX2Ekj4tnkoG
w6n/8Jaz3OZEeNqaCuGFDxtv9e5B4hoTho8pj48aHRroC1pUTQMuPVJDuqW+gEL9CHN40KTQJqOF
ictXwLFSKuUZsPQ3Dowahp2i+7WMXIaZKaRz+yrC6uPs20u0xH9yuioqapWplLnUQiTxThwJC+Qd
pWMCKVG2lpoWtO1+nNlds4vmcN07jTzr/nvtIFJXhO6ttSWVVKSueoQXWNWy/WpX8Q2yrwy7RQou
HfTfeHAGABJnwodXzl9OGz+pMBDVY6INyXoCVbewuXZZn7B3UNjSXylPzdDje5BoobHbLyIpGLHH
1vsAoC2mmBzuPqW+u94t2YhWrZLcZbpuDe2ZNStbkXg/qnwryC7hVCnUJYTykRwv29m/aXtZLVhK
jCPq4SPaoghe7AmT5zKlLSNeVGkWNvcyQ6Ng7vLOM0Y4J+pW+deB/cR6pJG1P0rm6x9a+yoClcFC
7s5vOAXWQWgL9dpzkSIGH5NBaOzLTy0jJ4SjqvfCXHgDdAIOKPEkbduRk33LnA98ZW1X+luJOnng
NFN+ptiBpSzA7Xm1q+Gltypvc1Ygbf+wXi8zO1SGbMLNSthy9vRI7P6RY8qwXL+zne7I9w5e2qI5
6nkP3+6H2rdZaacdooYF7uSj997tlSVimT5vIK3x7TjB7OKUJCWkJB+iYcCFZycXdWJwWDw3YZ8s
YrZE80PWRTzbYkF7S15gvFbOe04BqY47uGILnuM/R8lJfR3jK2D/6CKnSF4iyqkE00wwbIMRBTk2
PaCiSMIC/RHbdGDLvMvzpC86f5DWyR/WdEg6YBBcvOmfLIeR50015f3imK/6IlYzjePUriRgwWDV
dAS8jPz27wLLPjIWmgM2SWyIxfxExlPyvjmbf9AwSiG5u/BTjSfv0f/xiJ80OIInx2mYW/x27Kk4
pdkAXHMEOHXlU3zvuu4RrN2GvJkJ/Pq4QTP+cMWFVbSFJlXErWylcWLQzboTO1Aaf48UKE9vsVDY
7hJEETj1PW0zZFQFU4b+jD/n60mPQ/cyWaybaxbnIz0hk07uXHIPyE/67FJUTzv4HLr3MNm00yaq
woc32Ht3kIQ8FqKiraAVIjCscPoPAED9PohIqnqTNW4szw+TnmEje9moEugclPeRvuqyo5rHVNVG
5PqpOpah/KLsXX/8UkPkvSNpBg16/DGRN9HdShRWYjxwMjwlukMGfeP2vxADQ7dVzDj8DfR9/c0P
mlFfpW5YLRxQb0z382bHfHB8ro0rmTQxE5XoIWckxa/Yc+H1nDkfUSci0tgKrZd3xHp6LUQJgRse
WOTdMRPsF4OEym4DhOBNbwQXkJ2LDMlqr4Uj3XCDRROMY7le1/brxM+JEyz0qspLs35kH6DdbAhI
+w9uGVhzKI0llSy4xUPU8OD60EzJolCIefX528r8MRPWQI0CFGwdo4ce7gTh6cxlWL5PtUwu+a8/
xfKVfAaveE6pYTYuPrdxbZyFRjVI9E4aTCxQtuU6lLuBkDgE0RB7CkZ+n3wO6Z6FCpi4OblDYq+m
6Jw2evOqSieIIJCoN6cgl+RSI0w6iBZr5ru6LwWqQKbUqTI+2RFNLWjd93Rjek1KXxthAnTrMcO+
ccD3vTdQgubxP9UqxvQdF0ls6t7wT4J+tiGqILjaJeGybGhBVSC7L852fH4BvitHaqV9BYX6iQ3E
5VpZ2T28QdSiT2OIFXxCLB/4/BjNJdMtrNzWr7CkL1qQdo4MROsO/VJ4rUfYQ6f8TDRFzCRQnlhG
6k+sPvQQJGtq2XoRN/owUNfi+hVrnYrgZ/NGSUKNfenljU8Ed1yM3YoLoacu8/UyAZ38eoEru1iE
WPAhewIhkaPjL4yMwre0W0XBeEomsN8tMydyEgi7V5hlQ6SPgtiyl3Rl3/3iICpYn9FCnslgR/ja
4pUJIDGYUg/Yz5BvqKBAHOvrt72A0+FpR9eIkhoDv3YTnc6ygrO4cwM5RkI2UDVqBfzfTmw75BX5
yyKKHWwlRpMJ28UInAbo2+LCm+kS5yq3kIeXa5WOZ+1U1dr9XmL6ex8GmO5Av3bs0jkkE/bq3JSc
K53REF5BwyOqoNyVTSFGmoNN0LCvQw8O71lwbg1IInSOfpTdbAK1PYLIPMbcYDq/I63cm+oGP3Wf
jgYI758R53m+Mjj/IyVv4cr6N3sNRM+iIphtAqyujxKtgaH09nxo4QyA/qsbJ83s5VHvqhAOzD5+
vZN5eMo20T+DdPbM7OWViiXn0nMhaLB0IbXuDHZJJqHPndB2nlZnjsG7QVEoyWrMQpyX7aLmW6AF
F2P2ogzAlyYAh/gwoEsJStIFZDHU0dcrELVptR5DSVXUkgaxVz2YmnYuydTemys+SXGhP+Ns5bvw
OjpUGmIj8xWyWCjFByaThMdLjwOGcMnAKWk0cFYlsaH0okiE1+wk1rpO2KpobWbKLPOORFmnTUMJ
XQR/XJLrkLhxrSrwMBuz+pK7z+ORG/afhYjTKjhyY4w8UIwNgZmhCngfDLrYCSj99wVojKwmX9X2
v5PPa64QSVs1JXzuI0TxFGBIs1TOtE+T9uBcaHcXKCcejHiVo1YTjZWof3Ipxt9DPJorQmlHd2qT
wQpVas3X2mVBHMHKuGRvLSeU3laMMau+w8O/UUlpQvdRT3auqVwn22Ol/voFFXkHfrbT6Cn/GCd7
HuxCebMoM+mKCdV2VLlAAUsd7uO5KFQCJYgE6QduOrV/HNZSMFFBSti31UY/S97DccPyUHMSAQpf
Yy0DqRHC11nucKxAEtDaP4Q+1jOTWlKqJnuOiB2dwKtEwQ3qp36qqLa1CWc23uJf479k3TOa7S6y
G1KzHNcmA66JcD95xCH5pONv9FL2czw3JZPiLcFcg7MIkQlmQ3kj+fOycGewnRGsyAfg1jNPj1HS
UlDpv1zXpxtQ34lU0W/ixi4bu8BARF6YDk8kZFrI0N9jNM2b5Xj4Z6Lttl/k1TcOdXEBl752s/kS
EIeFDmThK4Imj3yWS8uZ8GWvisWiLpHzNfVV3o+CAirxTpicW4EzmNNh3Cqqiy32mVHl743hR1ah
zQw9k+TkTv09oJyukFeoj1xOcIUjD4AGNmcE6vpQC/6cHlKbRSiA29MkdpggmWq2p4Hfvbycjc06
UMM85OSvPwPhVRrqFJ641hCI4NV93ADqMNzSYdono/BIR8x2Ha8JnF8EfBJUZd527Zc/jhtYPQyg
iUJXCRSeQybXXsoACIZvhw7TTfTm8OyE9D4sXH658ZUiPiz5zTunQBmz2Mw3xfBmUqmltB1meVoR
T44I/yKgmYkjOEuowO18k2kFzPuAJ5F9ZHTkxrLNxcbVvhGRy+GLTybID3C6vJf2SFMRnUgVXjfo
f7FJCS4LAkee/CEIEQ7xg2nW93MLxaNkBcYk9GN2r810LKkHSgNAoEZNesgup1C4JYJXqneFYtOv
2dNyn0s+NyUkJx3MJUoQF70YZCwS2wzxrMjxLqd2Bfy7Cmal7WZE8dTl7Iaa5YhU86pjWa42BKql
GvcXG1+J7l6W7RmQ3WvDk6j5tFx/nwoTPbVxjt65MYQO2hQm93a23VpPsgFTrs9EA2vCuP23nsYi
5rgeCExz0QRAPMP1y4k7w3FI1pcYbO+uznI29+6tr3v5+efomwQ9TyS43xDaVAx915I4z+eqKgZF
m+BgaFhTSJ7eKOARx5ikdmWOTjDxjXS2pbafBE7q7a93slsf9ERQTY1YsiJFZLwbl5O16DTL93cR
++u1Gkm3DaZxnrgDLhxPEcWMEvMSR378gkH0Nbc4lVRXsUvSSY8xGGz1Od6W5M4Q3c12USRz5O64
9W9+o61MJmRRSETiIdFgOodHBnA7ADTOX7y1OERn3wu4uL6/jRDw7t07sG5P3uMFQ7+R/M+LNYOb
cZVRDi0KWzY1kwJLdyE9kCv4En2qVbuJhHxUZXZ3EyE6kFwFh4wOS4o7vu3lW0q/DiegJeoaH8uB
CeyYpQ0QS2iX6mQEe6WawuNRCGploUyEqNRRmQiKNZ2KKux7iocWYVqTgaRIJkPg8VZawSkOQHK7
cZD2Da9sDsawxgWn9RqjieuCOuKf9vecEdhlodDf4rXDLY/Dzkl7p45ph52i96hRI5hLdV6trL+m
8CxhiSju4x19HLjPkfzqH1MjI/sjc1II+MA7HdgKNwYwq/5QAYsLL5wwtJiCobRc0QoR4Nlb4Vae
xXn+AzT0K3VFreA23bQ+uIqJ2JQJPasTG+7Kc4GH7fG/x0vFFpJbt+Cn6tiQZip93xDHUaRJouFu
ahvQFozcU5RKnNfpDn2MIbLFY8s5qbsS5gMxXOdJviru9bvxrUfzqnoqDpTBz/l90ESaZnFL57A+
i/sZA35SEqJEnYBQGzUq58cRCMDAku6ClpoRwxPTwpE8OGfB6FapuDY4Z7UwuULf8utiqkcLFljr
SpyGUAIexBhJYmKx7eDWflPFJsDVSK3HGQEqARfIsq6Q1o5a6reeSNKkpufsEg8hgtiwePk5XmcL
qQ1XM0GLOo9Nyux1ew/2mSLEA9TFr+vYbES2lCoy/lC6rLXizbd2sZkEt9enOpku1ukCTCrW0c+a
NK7CAL9YLol/qgGMOGFSeB4GeV4j5XjRYctBoV43dQH+4k1fWSZ/p7ZHIaS7Lj+O1ZRQtH2DI9gx
UHKJdyiaU114wO+fx5N1U24ybjlGQvCWlVdGZ6qOMOjDjwgLQSrzuY23HDidIcFxZgBPlEqHdgrS
QzLIBYt4hxRuahjYnL+QfacvL/QYBEgnVG1O2YoWBvmksuiS7V6s2QaIb+0wDi9VA/mMJdlABx98
FUNcEnWGABiBJzx4rH0uqOAYlZXtDPfMvcdd2UN5vcx8rbWsd10Jnoz1hfBUG5IUV9nLMTx1JrdS
AZXAxJIE1kvVOw45hUvgayq9ve9byCPfje51JXqFlkmIawS6Bh0d0/eeQJ+Dh2SmKUtGsJjDkPWl
H7mKn2jIXhRdpqLvN6J7AkH6ROVf+YwLLoVHRuCMN4uXw5hMBmrWucsIzwPTIAb0jx9v3DPSnuvb
kSrAMPVUIL1pPS4tpT+cNlZ4eYs/HXwA6xqj7A27e/B7Eym00dxSsH0kfEjlEEpDQFcYdhbQxLUq
1mqEhvseVJrvU/Rk2+0fhYTu4hvuenD64xHREW03s+GqPRNTxp/1qAeq4ATpVSbQKOgxj8t2NkjU
s+fzijPW6kb3BW7eaXkl841AAlPtAc/ClPjBU537bI0gsUlgVO/pQglHl9fJFFo8F0daBKV7YI1c
fv/c2IS2Hl4uzDI0/UWvw9TUaJWJD7R8wcGbyHY3IpGmqoL39qa3QVTD15EYkJUZzhhxcK9TgsdT
rH38lx14P19+1JbuJ85sDjRdgs6igdRI5tJHYi+EgJPLq5RKzPSywatcdFvYOBMcGwDY9jMpAGYX
AHRm142pf8J5uG3w+j2k3mYtuw1qCGsIxPzP+8vb0V9AbzcSTBjBaRXQTgfgxvRG3tOmiJsosqMq
Go3NqmCdStpVkY9eQTL34rjqnm68zCqFVwPbjouPVgKi4kCx2EdstRcWJRmY2RMN04qClPXJ9j5O
/w6pGaVEB7je3wF8Nxj2LXRjC5UUq5JCOQRNd95H9tnYQUNQDQ1Voj/LosbPwDtHZmUMTas5Z5w2
IBcvGXGTht7KPDKireWjuEjqwAxxp+FgH05uyqPdi5GkATy+iwLeRfErpzsgyAsmc3ILsBBxIUWE
2VWilE6Yw3zSzkvyIOoJwGUq/81/jkrbh8bEMyD7f/ee6bQd1Kt5hKR67NYAaKsvN3MEPKtApNJw
RNtTPyktsTuKpMWJeBfDdVUSDr5SD63yINvsz+jxw9ZqtPcTwKwdh5v7zaw5U1tOCC4cEgDypqix
pvLnh+YKX8GpR0om3TrCLc+T/KZH/VG9+dykXiFwcSISN5DlBWA/rV+fNJ+earY5KA+7lhzHqz44
CDYtu4mlnD5NBpLO/ZW3VbD/DyXUOHs9D42Ja9GwFKArPzqDH9ufRMwu1FVMwd9IrmvX/kPWdCnC
bJl9FW5jXpiz3E7ieArVRHvTqlVKd3HRzOzjgjsSYLBxqgP2Q+m7e+Mz3cETS3QJJV0R+NI29BjF
rm/1fObQeTZyZ6xxw05vgI46VbLjlNWslLF1TPEvmt5H45VbIprKSl4KbdgRhkG6j8I1dJep1Dv1
96NsEeYGW+oz1BsNESrkGZ7ydWKIZayO05Rodkvo9c8aJv9OnbA5Ps8uDkLKEEjex6SiJB6FjKiM
RkQ9KnUfdfax8MeaUnkMV7qonWCJ5BujFHi6SVmO3yTd3kjMgmGOIgwogZx5tFN79LvyjTrvbIfl
YJclFyOglhH3I56zk3jIfsFBRtCW2sZE2cpH+Um3EaQ0PH1KO9G+x/7gYGu1efi2qXWaYPVm0OEU
LA545swqv2GjabiDqszb9tfXKWgs7fauUSiUphClwpg8WKoQXEmsxJrkVDp0HDOoylZ8hvCcklUr
K6ua2VGYD3JPZuJ24lNu3hPVm3WjYgEqtxj2dmG2yyRyCajexFO3HxfX3RYvrnJb761jXFGYJaMD
NbhIpWRcrL4AVmN+uB60POwHOuYsFVKAAYkj7qA2yySdeIpztL6lYVADza3qUhWYCYikJmKE5SRy
TxOs3wYP48MUtlfXtXvEREOXajNbq4Bui8hfHlPlHl3N2P/Adb/gV5wu7pgMrW4OT/e7dTCcV05i
jSNozsZ217O/lxju2j2xmlE1pwMLgDut6gP3bv8mxsZj1MZjYIXXuB+YFwEtV84kz3eKcaIq63Ju
5jQluQ2SbpyG7phCOy1RxGe2i8X85oQot6pP187M53YqC+zRwAIKoOKEho7VtZbQIv6vKKzv8AtX
Biro52vyy7UtQegdUewSfXSjuSyqy4Xuv5Ex5SiFdnPWUujDnGW8ufReTryZZeZa3WVi/yWROgVH
1vfBcXCWRUO+i/ubYpFChbHseK0nH1JqJ5kDnYNfCW3XTAsFaYGa+e2K4cVN5A9werWaP4yuf7vt
q9lkjHqPHw4jnyMjtfgcgWDlXEMXYVh4aPXy7tk76vVx98c+L/IOPfvYLktGNLPmxMvwjdyaA6Qw
/q5WpSjHSKdtcrr/Yi/CHvk3FnghG2SUMUh+wurBRqrWbArRKE9eEgdJUd2adQI9YwMnuftyDr1o
m07iifJ7WOZ3yNtRnHGfX3bRjFvWhcVRIt002d6Xxs3DYN9L1VndWL6lrTiJ2e8JYEobqNzVpSrd
P8oLxgoE7os7kKa2TBNb00RbCHZL9L6E9IGZQE+XQrHS3S7YPDR9+Nenm0Gb3mQdM0WjLgOLiraA
tjnbgu2z5+RoDBtq9PGmaYpT6GxbWR1PQP55vbLj0Uuw7EyeDKsOKcP07Dg+9ijMhvenUJOv3++1
e4WDplKPOcYKN4QLVBflOwRjQTcv+s636taL4rKF6nMj70iuCPHgBWMv8QxfPg3i9M4hIX2u21Nx
hhnZ0z3hsNj18A5uNvX4UymtUqdQg6LbDHnQC4uWAEU8lLZj/oR5vnTqgw1uiXA9VXuXmpbAfk97
fL9WvH+oy8QQlUyejxqnI5FOX92AMLZZBTgxn9KxgwpzI0uXyLcPDXaQLLCGhb45jNZD/ZyiemQt
mHSlyVZpYxygH5CnFDyK35c+axNeWLy9oX6QT8aQYwtSK/LJ9m9W6amo3A+gqtZIiSmEW0zPu7Sg
6Z7mBxbu3MZsNq/cjWY4MJRVg6mLr0JZb9PEGXusBnvZ/7ZJhCpDDSCv6dqz62R3Ew+rpFZAqap4
5CDus0yNIxOBmKOXVxI7qwmInzqkOcNBU59bQQi+6xmWDurUeNN6vux/WWBgbTPeA/rB7uKwg5RT
5cLqbsg0HKovQCeu24gn84dNC7fygAnF2oBFhQ0SEG4b1V5X1rxA70VGCFHcmrxeVas1v4fnmg6O
EgTHXubypQNx5AuZ63NboNBxU/MkG4jZznNpcHVdiFD2AsTpVOgprNKFXbhUQRr2nCADJXirALse
FcqRlbC1cIqwggSTd/Af4+l790NsGBgdweU9Du3NXErik3shsOOEMSE41TtSHep8Tw4X21kYvUgD
8w3dBgjg1Nr8dYV09gy1EOvscBZUqx2Cmun8pQIK6rUXQxZnAf89FOpwcH3wATHxHLdT67ivF/Wd
4A//fLWhYJuWl7SHew9C5VLcc5UL++ZLhYEMZtVahESsNYBBAodZu0dRY/GWvuIPPWMdyj8BtFYo
SsP3pJm3s5zbhnWx+KnjsUYMOHJ58e+Tx3FkrBhitcC0A0rlh0y4dswe7ZE7cgTHqi7Bkwzv5+25
Y0TTVzGFTDmXl+mpG4vDKat8ZnkfntCqAlhjOc1AFk1A5jXoxTHSKsMp6Sv/Y0kBl+wC0tnlY2e6
8eUYxp5DEDFD2Gfw4G6JmT9bOCgR6ScMILm2kw3GIrr5f5PQW/mtRDfvN4lO5BGUVwAjjKUxp6vu
q8mfwoCSUBfL1nylSz1KwrC89mqce0bc9bKeEtVeVuRKxNpTNp4r7MGQeVBjLe5xRGxEWQgb8TJ3
eSrl85anGaNOFbxhPfCBBHb7oaU+XnRbSLNnCkWQ5NJKS5jRcNWdsmqd+TQ/WfYH/1v74QZfsUHE
hUHbbMsiwvj6Gs/R+COPhbTTj18cwEfKzvWXULK3lnF7PSNd1a51JUv58bGJHPz2solgP0cG3YVC
0AAYP3C3BMbCPi0URQ8fNSu9yP7TqcPTGguDbIa1ND7RZs0JWIAAvH9FgNxbMsc6iOh7Tq6LOxlJ
OefdzZ1l8Q/hu8FgIhBoaXNptYg5dIF0i14XGw+LhSEeb5aPu9Q92pK3W6ttZKFMJbHvzYFUW+m9
MjsJn3c1LdgtAkAj5I+UQikJyC2YNHC2Tkt7xMMhLH+bMZFkfUizI9+Txi7EwzoPZXtHlw+CbjSf
gLqJMo//bHljaMpsjso1tqVDB/TLT7t0PiXZbr/+1Ux55+ee5QEFgLSj0smqdsK0/YDRnAqK1QDK
owqxVNXI6N/ap3O/uhjXPivvINrYs9zqkwYubolnETqtSnI6QM21QbrIdKjXaPVKyXHYc/2YUe8g
BMiCuEyf5ooKE0QPQltKzoT3+LEEoAakDA2Nc4rqDulN3cSIA9HvYtzevM6hcLeLlDSV9koeWS5g
IlVJDjSmvaGPAey3Wc/3dAJbFryKdm6LUXVZoKiBqx5nFfUjwKk7qNcOHQjNBR+lXwW0Eu772aB/
c3gseW/R6qKJtmuPoHb/1TR2qyTTMKCaxV96t0pIyvWj0yTbVTuOlQeWsCHoq8UZ4bhjfG9GSmhQ
j7JbsuRQfI+/JBSlSRjO5GRIgDJNZ/9X91gHfXWwy2hrwN7p76Zt80qrPo/ByEAtvVaUG0jPm1vV
Z2SoQVdUJCSQaMvbOXJw0vy/i+tNnbWUHJa9GjVTNmWcKY2LXvf7sfGNa8YN4Rsy1OPm7YeEeUy5
V3LXl6+YDxmezpI1WCifrzhPz2RnL0PFh0ZnndV1B1EC+JavmX8K9UIvYvvN1uWq2v5Z820gjCno
1qWQ8fIXxo2jFm93kHOPQhSYBsB8Iz8jIt0B3O+y4jo/SD4skc/HEKLjB9oUFWQHCqPXHe7cqHtA
o+T7YYgg+0he8AMHykmRIxO1wrIy0EVf2TShyxf0ClxstjyMeWOfmTLJflrUe0pnX+ywOSY4uJiB
uLkLPqrkEUH/++Wt6NV/6MbKqKA1II4UyE8K+4zrXYNYUFDEd4ddmVoHyRzuurCi5JetGCfag8gl
Xho+0a41JYqYkmSbvqjkkKzKh84GOrJIalME0TxPGX/+PRKAqepXDO057IIe0X4Isv/emlWIFuWa
NFBT4YtfHFVoEuBpSVL2JGKMNYqSegq7JgMbNseqF1oiZYyQJez7NYnion1zJR/vr7gy2XvIi9qj
lppZoxmdymVds2vQhdbZ6o/1zzGamrxKKOX2Z6aqanerGmRGjnuFtkAX7G0orwMmUiCGevYDiys2
JzjclqRq6r5zbRQuTdj8JvQXTqbaoOdkT4k5sovFOlS9zPOFZrZxg1MwCVrt20kbeTg9kyraUTU9
jUb6P95Mft3cBQTVbLBNY66uOY3nMuay5PEBLa4CkDkWu4YO89TdhOBrh2b+1OsCOS9gQYfS9gt0
/KnZ0tyoO9sh3jAJTsK8/xdfkyZYiVw/okiQHiT8max2uWv2XVZKq7+/Xbm+epzX4WbgEP1h9AHy
xsdcXMfL19kKBu0xYmlNBtc6xdNxosp+TubzVviRO2V+vA9n4uKcP5vOkXMhfVmKMtJ8YqKSwLqt
CMYT0I89sclGPcnldBjykpwDpX6HYS0nX1XiqjTeiq14grYSiuPSP+pfU6Eo6OIuDCq991wXZsZk
/uhflGrNOK56aI0j85hhkFUUcWZMNTxS3Fa8cUTipJyGgJrKOkMrKgxQQHONWM66QaXGMcLNxBT6
4pmdNuaTyxg5GOaSFftuZBP5ptxaoCyO69NnvfWRsvq8530R0qOqxTA6lUHjqwt2fK6vWrmWrnkB
NRynU4HkVp5xbGW8nTrLpceMNL+ck5twfRKqrVp853wBf0bb3FJbvcmvwvmSk2bu2SzrTmTsV0WB
LCep0vIGSKHcBZeekpTCN4ck1/CZofw2DLMpGcz2fPsWjzr5YVVnrp/Gw9xz/kmA//8+M+V32dH4
Z0HAwFFV5xQXdmj+c6n8ZnTT+57vqC3tuw5X75TpO7Xby5ewGyCPMLqjIyE6bIHv9vfS7JztCYU3
8Oci1qyRbWsA7udLpZqqccZcjbP+XsM0a/eu2WbTR0lzJe2knqfdvXfgj8rXJKCPFeI7Dd1R84qU
WvVBNjPs3/WxMLi5CcQs65sR48cvXxA7v21BlM9cZkAVOEKj1O/tsxqmP0iija803H/MXCfyX1gR
bu23rjtbBiWA92Kda2mJw7faLTrFICz68RCVqFhI/dT+llBthpkMPAlUvYMNoWD3Th/Wfr+UaaAQ
77x3YfYrLxcXd2AnJ/pdnx1bk1ZoJ626x4iDMyPUM5h50sGUfopnLyva4Lkx7ccU6H0T55BU0EQc
ojVyRsg9QVqOyJPuTJo8yvs8Zm3l3BK3E6ARJH1I7eZ/lGDpESnoMM4NeRqQ7Dhomkfkw1/SnfqL
QVuJaBHtGFVotF2MHpKgTO7I94yWEgfV7GwZsosHjzdLg+HrmJlVHwoo1Kgk1USWuJ+8WDXcbFtF
9yooMV6x+/acl00g1dfJqlSgnKzHQFpNjJB1V3qKKwHVCgPR6Xouq92dd2Lh6cAzTHxVsZD+yYX4
2gCLLO3AFV9PO3WBS7K+PJ3e8atyaNtEelcAZ/Go7FkZHsKJor4kxAfJaC39+of0eQos3tVex3ZM
S0HPF/S6COI5/NADmJyDypnr2ZnI6nArafk5fkt3z8Ot3L61k7hdpzlQFwV1VwFN+GIhjhBWnoSA
MzG94GlShlBzJKk+/OdoRc53CY3QNr6XZbMDbYmJzITgR3vobMnUI2s6wbVkm7eaL1eF7sZnZ7y9
TzEElJcbzRrJ58KapTQgRUck0Ak/B+Z81HRn3WKDQRRRyZyX5BovBY/Y/z409sUQKV9mfHOl0CvF
62fAMr9l8gwkgRSifA0jV/8Pda2nEmn+aoYhgzYrRuF1HfHwkXpS/NnQXMZP+6gbySormho7vZgr
J3fH+K0pJD8XB7NzGGOcdnltQrDpGUsfzWRlQJ8ohQQU2SXo3PIofYe6AV0dXhOPDY6zuUbhrayM
52YwD5DFmI7BK2yEZfJH+hmxag67xHcEKtmwYPKPwzexifebSz8AcvYBGvebJ/y/d/CM2OpXKxJo
G/dz5bW/eMFeeaxnCRCJaFMprldypHsqm4XAJeZhQOun/8YqhO4TBVMA9dn2ggPXAvFpyvqUnrHe
eFWWzvddZilFniG1tANOzVp9fPiWE2r4jLnctnqU6d6MnilHSTi0MAG/K6lLTBuBWkkt8bGRykjw
a+ZmpPKHmcTWM6f2ttJxfUGDktsjo+HYkFLUp5pzzasUs3BGiI37vN79o96IWBz4VrNdhXNDoCMk
+M/xe/UR6kPAO/XnB0cfKRl9I0FYavYm0gy7XAjp3Ok+LBNfOIyzAJ/yr0OIKOiV07nBth37jaC2
wDXBJ1wrfVEsaMbpP/93DZbOxZ+wOv/xusa145pSl9Qg21l3zsNlJKABsOE+LaRajwMtyu4r4jF2
rjA42QGy0/k6Bz4q1c1IGnASjE+hifc1vrcf3Xvq3yamQlxCx1YJP/3ZpJxUg3OjUM5t8L6txAEG
YKr3esCVbGYHYWZsGtcejaVHI5POdu4ThmbC9aSSCpkeuSqQZxO95ovWzpJmznUwjw7sX0WTOIyW
h30UXEo07OwCdWwNxRRxTKcNi2BFm7m/jNJp6XmxMrQfsSwYOxVr9Q9aUmwXfUb2DfV/3+B0yAF+
Gh0wAg+e68+Vv8h0XvUBkttAxTBEW73R33oC1gKuXq679KeWT4B9D5GMEM6yO91SFvYef06QN7HT
pCjBF1TONZCqol/cL2hTg/VTjYrIMnR/EOoftUZOnQXFgRYxAzLMQrIAUCtWaRw8lHlhu5C8XC1P
HgcpDtplBSaj5m5G8ugB2vKcxyuyZbYnXfisZ7VSW42c1s/zeLqV/50VNBs06OEmq3Vyk8fK30w/
84jhmojv4dPUquOThby/ZA5UcC5L0p/xIsMsBFQBU1/nxX76zpGKmxOIK9VNp5p7EQcyxMeseZpV
bSyTaGALNfxe+gEUEDPLlxBcavneLJrfvnButdSmPwI2QB8YN89rRTk9TZoRJLRvYECIrGu9rp+2
BhsgxWEK9/4FhhTGygEQthHsWsHFHC1dSq+AqY4DqkPeEYfOrgiC6pMO/SZL0X6iABRdyrac2Xdp
OVX+a6kyV2s+v2T1XyQqC0XneplbK37tV/9nkpovYQp7B6pJ7TU6Nz7+T2vgoTbL5QcdQgrnhHwy
tjSHjaBm4pWZsTrN8jyYBfQdBCoG+DD9HHb5OFXQk1V3YStekxmgAyZxX5UwXi5PjZw3IybjtkEf
0gHAbGIDSJggqoaYLBw4HtcdBJxrdh1v7/y4g6DoApJGyuTpQnkK3D6CUnPLYi5STXPRlpuAY1UU
/Zpq63MpngBrYPNFbAKuzThDmwVk42Iu2B3XfVnaeLtqqstDsdKlA0BClcM+iBu87rdtF2rjBRb6
kL5BC19kY8caY5qGUBE1vIUYpHHzbodtI56NzrxmnrWuXcVHxPFtei458ZXg8S/klOirmd7qBUYn
pe/Zq2tqSxAE5ZjVBXw+PwR2oq3sjEFm1GjoYltomI+Qq+JnNY7xODQFWoneevsCFbvgemNV5KFF
QvvdWp4fNd2CSwVEEO4gZF6XOgslSfp6A43fvfTqe0luQO7Gf85KfSNIeYM0O1t/sQgeoHJXVYAG
BTbL6bIeixHslzLa1hmYWrZfEUeD2FrJh5YV2Zr0HfCYK5I4G3onBnEDpKYj8xtG5F8tyLgj3ys7
O+NfetcoCOsv0iy3pQE8iiMFVBflbgvZwRICMmKNOiL0QBomsRUttKLESvZGTD4/n/yO7v8hN1OZ
eI4ASs8nsJlSQm/A7lpdvzClORklWoVSTS/U1CzoJnVV4VrcwAbGejMuHuOwRmcA6FDRhyoMCRKy
JCl3/KCKLwrb+DssMzkUbkYhcS/hjlI7vNw+VK9A1DEEdNz8A5bLoxN+ig3Ga8rLou7Yy+63RFOT
YhvpJeCxHfP7ODRjSKWrizdhcPo8dPrZF8BfViujzJkT1BDBgMMX2Isz+1WoP5y5+wmWt80Q3wac
xUtqFJ5ybAgXRkHzAUqH2TkXLY5CFb9CBTlNHVcLT9XQ78MEpRaDErTxCXKkUX6SwOPBB71cnopZ
EFGqd/RIVcilD3QVoeiXTf4v/9812QuEnkWK2fLU2pCmTn2VPqHuYmAr1WTVPzn0KHzjdEfKjDBP
SVrqcZ3EyP9szbSgDHZOwucUWhnCG8gY5O3kQzOCqKUng5D9SieL/OqWsjT29Iz11ZuZooT6zK+j
QvrwcbJL7FECIiNcKgI0YP4QjFzTFcXhX9a8U6hgayQJ4TGCcfrSsByAbcm0MZLz41IlEIvkgfSr
IlnYy3hJYzO2sqHFBS/71pPqapKKNhgJhzcgAWlEQ1GfshZD9U9JOW2b6fTu0CNUy2WYG9Db9z0x
SUGZA1DwgxbOnYp4fmYcctY9sh/Hpht0QH/4U4Y8Quo+I++BAlmYiS2NAkliheDTtODlj7tfNTzw
ffY0QqelNkq2luYpFiyGt95+AABmibZ3XWXKIRsv8y3a+sMHNMvvaT1JypSmdoVTSWuE4ldQmmHF
QU3D6LDwxrDqBb6d2gRqBtRe5wueFnwhciJs9hOp6CPWwmvT0uDZlt9qsFMEVxkqcCL/7aAo5/Xd
qRvj+2PEYIv26/Ff439qFaA5+8mO0yCi0oiSjglMw8wTHd3lH1GzmU+jCuERkwiTU0DCtB3lUIWE
YBjOdIuZshLDtrU0sv0Fn7W2vCVEz5Qi7mmV5nFCtR9js5t9+hSHQoy1OyV21KjfwZ8+vkeoTTSK
K4T7xagJItq00aJ6NSkC+6r+2Fn6evdC9VDZ6HcZlkrxT6cuFOWgEghIcNhw0B0RONfI0zvBxfHI
Byc9J8gZfmhb+jAUrsoVbHlONHgKzhNs6EEMHyf+Xwjtq2DeDjWHiyfbz9SWT91YDlfFt8yqN1oB
knX2xgseU5MDyHMUbHOlgeX85XToFLJcd7YYJyG2mwBDesANqFeyFFnuwgQWOBLxPJpbG+u24PVd
Tep7K9V7xubuSIGrehHmUqB4A8zHaI7Fb0fsWaBLUlPCriSaLpaRIlU/oQBlVdDyvldDHMgR/G/o
3wbCOZzDbAoxLEmWenDlYRfInwRTtcQMDf/YWt+0OhsrBoo36mXvLtRCe4hwQRIuY7X76j7fqXWg
esCI3p7sM8Dy58+3wtWRlO0QMe4Ypye7ICjK1fMH/JhaJswp6eaYxYN9pz0RXbdhXJ98Wp2DIf5f
HM9Z6sx1b8XkZjxMF6skS2RwFSFFHckKDv1M9Zns86qbz3ftYFKTypZgKuRcGkgY6W3hA3cEjD2Z
QAwxKUfoeFIIv6ELYtW5zdgXpLx1DMlbLFkDALI7hZMhqwGLlSght5ibG1yGT4zImLx22PkZThJ3
9zOXJ3+kGcJfHDLtUCYbHX5KwKr/XJOqI391xiwebRdEea6TQEEigS19hA+C1b8AwBn2EXorP8fo
vUVhizQub2rPOn2+BSCkh+Wm91gjGmotmoQy4HnZ59U0DXTGJpClJztRQkUvVkbDvsvlmqiWGIEO
cs2GnyjLmjbKGZ/LkE5UHB3H2NmIqbue8BsiplGVULBnTxaWGxv26bOsjKzob8ftL9n8NP3q1OBn
uHO8i6U+il9v/N8DmOoKHlZwbAH5VLT6qniXv09smhRyR+ipZqa7OZjKogzPnO5BYzIZr/HCmNc7
z795iNG5YLGq1x6UvlwhvYEPNfZSv0AKf6CZVPU1L+UsUhy1fAvduawwkngobIOjKZNcBLwMwBOP
IXL0nQnWoxxRioqyTHD0/SvBq4RaQa95nssMhF0uGcvNboY3WHIPq5094EVm7YRa84+/7tUec6/L
2Wj33ETMiry+bQY9TUJ3vHegrPITmdEqXwusD3i64fSU+xC9dwyY+BOXIRQXVCIUVmbrypqGLMII
UAVVfnXuaMIfnBgxW5RFK8yzxi2NWA/pjsi0UB+lTEsQdh+y+zob81+J/Hh7WSKWOPv/+6jasF9c
wjWrUyOL9mw3kDuN+pg+kX9trc+UUZmRTrnkNWsUNmhL9l88qKTKZrQMiDPjNPm6Sj6xz6IQPp+K
dBGhVtpGJT4UBMXIvL4YBx9NFTWJORRE6QcoVzTKP8zN73KeXnqiEoBCueS7TRrHrf6DZmJdyEGh
llcBpKlpogFmXKAs7ude0ls/IfTg9EwkEnPugkkXF8akmwO+S1BEHOufpw3Xlh+tuxAGV7rPa+gD
wClmZwIJ/D5y51D0PxBqum1aO495zRFi+x10IHuxYX2LiNUmwv4Qyne56kzLEgXROhb9fhtGfyJ/
nnz25uOUDIxskqYC5hiDiOPvp78B+e7qMkAerPjupWmdUCgHLDC4hVjU+KZHLRB4rQ4veZkPsX/c
5FQMy10eP7H9Gou5ZNH4vqzYDfSui0tZMDMv6G4W6+ZPzuka84tik009FB/2iTKiJwURCXJw9NiE
ReHKTXae+GqCLCOyCEpWNrctaO1aefYgO18/yJbJ57JO26Fwll30fQp5by/O/vtaDVeW3SvsSGzD
YJGFnXa5Z5LSTtR/rx9cyEl7ugDBtbO4RvY7TJ6M4FXc6Rp84R7aFmW5xCU/eXQ6WzoZvB2Ml3Kv
DgFSvzNWr3NR9dLYlpM63hjbWw/aZsqshxbhrCWnPW2HlFKZGftfUF8FajoBk0/gvxohLe4zGhyZ
irR95+OHiZPD8dDNiBuReonRT2wKJ+jUzjDtW2Nk4DCamTsBPpk3uetWFE0GX3m4/jx+eOYc8Hj1
vTHT4Mb8O1cc61JyDtpYXAbAKSoKEzsr/VG0jKig+qmEJMpKgwlKXXleKC3O6eZdYjokinff1Eyn
4xlSBSlOaGUObZmnWoB+2qbp6ZmHyaAP5umvcxCa4dcbB0lcIr8hPF7YpFmrxhWwRPPtNs5MqbGF
Dxqaw/vpWYpuFjnQLpM06mn8+S3/qd+d+n0YIWy7hF7kbZh6yCzIKuaAigerY4BaVyJksNCJSupk
lurIRL6m/Al/HBIduoBN+qpOYcClLX6C99GVFjseHBFzCheZy4K3sTU8RJ1/rmNL1FZZ5LlJykZV
Jj0WXtsifXsX+yYP5hmZfHQMMemw6DyEVOQVr6FWeglS6I7VoEW2um6OJOi9raStcXV4w5LbfmoD
d8uGaR1/kzHuss9qwCw3VJNMNzBRTSRTry5TcAkuecKGwqBDvBnt+KKrS9Mn5hL5ap4a7Wz/GXPD
gcmOg1mcQFoDwAOhOewMPiRABzbJ7kAG4WOvgF2S++3l6CdBF6WBsnfpb6nJXkwbbQtF4vIjIL0E
ExCZKlY7I2SXJbyqYqYBUncBF3otDA5bG4IxIBHEnzLteiPqCLfkc7quG/h6WJKox5VhlTqVYsjt
HMP4VPPoBImILbv70UVrX3/MOE8tySo4SurL/8GzXuVpmwraD1TRazY+OHnBaY0wEz4voxAm4BGI
b9kyD8SO4Nk2Xqh7RK+ndw64OVk4NRlNpopyXcfCz14l28YlLRD9m5ntui06nBRL233pZ1ao1Nh+
00Yeaqlon0otnXgdcEHVKihu+HjjpebcgyeSAVgivD9ShJdxZYnYTPNkIlpCiRbjJHIxorPbn+6X
NPosFOf/KVvB7jugzOdn0XZczWO+tUdmbe+M9TxOw37bZ7bJMvFP86nzZ118ukwYNSGbUkHuXMea
v31Vgh2Da19ObIwyXbnkgLzBzFMhVHiJ5/23g/zmsjH9mshU1WFWfT8F3tjUK6fCRJuqv9M58tj6
mtmphQw2x9a4rFVYuFTLZHy/6xmmHs+vuxbZLVftjtLOETcq5ORy7CmmrRaS/RVzoQ6kkaRrpmW3
MTXIbhUg5SErPEtCK1ewrkTKCYAshHqRDkdOC4hoI52mvo1kiLxWznKoZY8zPDgieAiZgQha1eW5
3pRvzLFvgCZT8IOU7ToJwtIXtzxZ9PDc8rTukH1gGo2NJSJCC8dOANbCchCwky2y/QqHOB1/Qb+I
b+bhm9FoHEhU2m8QDRNqpbD557Yyd1RiqVqa5r4w2/BNru29MOcdhAEJc3GjWdQJdls5hsW4c/5w
K63ZKwhMDuc/4LCD9HfKPW2NPI3wbcui5qz61vR7P+8StlB5sXmIu3uIH0ZAkpswXRjn5wKsJ6tF
/jiOOJL5N3VYX0nkfgbPnRTpOwDClMJpTXRQiOsdsB8v69FC/urhokvYqGlzi40mt6S7sPoW2SOB
iD9lYZElnj6T2nOaYDToI4w/tDrBJLzfDu3F39WZUidNxycsDORLydXiOyZdIRvLh/EQO9p3yxSR
hZzWUWispuZ0muBPSekx94vzdf92Ogw+LXEcWnNKgr6k1ESqigBNgpJfjZBBAJNvoxWbedtid+yE
U8H5TiC8ZpDWTKa1skFJVhu9FDhPKLLlY0Gqcr3/CWrWYGBqHjigMy+A7cchWzSENy1xRyXvDWhO
Kr0kBHKQoo+2J4a9j2D/u8kSupHokpvViXcTZs5jb+cAb6A3rGGDyWmembSuED8OMpbLaswVGrNx
govUae968UgXLn72y06FM2Volv8yLpqmQSQWIGgNY6A9COgxZWUoipZmNwiZqQh2noXQfvAJEZCA
TMiqT+kzv6cFmAnD137zB00l1d90TUf7LYkmx/mDQpSe0Z/K23PVyX5DfaAJTi/wxUsYQOMnLB+k
YLu5mKqbKQHyXeTEWybxc7eEmEtDy7PVRu6GtZwzf9LYKeNpfjlC2NIZD6wrfbNOC3/AjUhCs5Jx
a0WGdK/5qo/V1ViPS/MkfB7wd0SV4fmKbtYDodDLTTNz/7hDDwfB+1lIA5k22x25C7Hsh/bbSv0C
X9Wu1BP3TrIYK2AO8bcxwpx0G9Z2w98JP404RaRDgo98alYPhbUkMcA7jXeIRgPkZvBEWk6Myifm
UYnRWQo66df3soDiCKoXo8/2BuEqcFKMOgTRrjYDgfoDfA/oZfnxiNi/eabRMYyL/VvuRQpT0JrY
sJCpbI3uTamu25rXzeEaGRk9gdebqGujW1Fw2wH45bWcFdKPX6rTzHelQGGydUcJo7k1SSSsrehQ
gfs+tbokk+6agFhnU0asA0L5tgiABjQZBmKnVIkypMYHIlNHSw/Y5+3UkRResI0lGvYUUI+lmimQ
ICyzvkP6puJca32RxjWz9NJF4jzoOi3Xj+zN0HHZLRwPCJZrdHTadEMF84sWhU6HoGyDPFXZoRGu
FTUEujYlDAwyYO+Mr8Z/deagE4zCkk+s9iAW0MzMv+4kZaNt+UdyzM7Ijiu+/ObZfa8fBfgb+4Ad
HiKoy/AhJi0J+KhhyUxbWCzk4P9TSO2/U/GAKrvL1XqWAR10DX8RXFGhyLSop2L0nKTCnpl+Byc1
XF2weC1VHR0pvk31DJzRxkqlmzPi6jw+sN2RBsbzoLDfk+pYBIoFKdlBSAHm2m0sUH0n+bQVuUHP
jzsL1c2HQ9aI8gLyAJOXHRe5zmiSGPg+o0kFoComuoy1CP7py+W+acetmsRed6waNA/WXyMHG7NR
TCPP6vTPvh4mp90FHubtRwOxsqbZVV1DmEBE0d9jYbIRYC3YCUIGjhwGgQbBrAktI9PN33krcAZo
RwEBs4KduYjBW/L98kp5SOTUncW+J04Sz6wR5alQoGchAoGpF+/wa0XL5LRgAyET6ifg0NpLGSsY
X1sbaK++c3FRnH6qmPqIsxAVGHeLQykahFYi5AMpQK75vr48CadwI2fJcKWguV6OSqtHvzfgiZaE
uLG2AFOKLBSmEjdJtZ6A4j+z0Ahn6NU5hYIe4G9P3n/rvHuXV0ILPLXGD+PhU7DRJStOBglJnOYK
2Xibatrv7yo0COhNMpVQeXXkUWZINTq66UHXJIeXr4tFZYLwj52Ah/9p4hmtZMmQxurUX3IFZrio
5K19oZFEsPdDD+6ZI1EDMS3G8uMeILXJ0/UwzKbEvBS33KwPi8EtZXOg7INdmdZezcvF8NuW9g87
XsdKBE+vYlCQ4aMIIcNXOHUqBbbKpzRFm1cCqKb8Sb8yEc1ftJUNKRdWlxmqWmO010Hz6m5AIeMK
Eiey4NdfdZ/jW0SzOE5UD+1ookSNKP4nZ+6OJCoEd6O8su00oV6bDmnZJogiPdl8e+Iw8Ea/3rl7
mAUI4695g/AIShNXGYryRAXZVXlYbe9+V2IJespO1QW1ROUO/sOuQC/Wi4MHHRQLbRCuOOzKNV9z
rzjwjK3u9c5VGgKGcyWU6/XvnqQnkr9/pUlM2v6fOCJM/0oefKKL23RiCZPf4XW9piGenMEZ1f2x
8MM/nRvxP8ZVuE6SuaW2d2+qUOMvAkPY7BZ3Wa6JgxQWdS1MvQrh/odqkfQb8n5krA7OKfyAal2q
YuUBAXpNlTz0xxN9SZaLqH2gx1YliMF8ExzIIDTzJy0pkJEm4Cg0X/LfDPN/jDNda2qSi5KRQZqV
n4J8yGoVFi5mrr0hnEs5zgflDooccyDzRa80uiZsQOfogfPVMJxmhJsrBCL/22m9ji+TMJGkikwX
7aiPj+w/TynWK0mV+RvlbBmy1kLLVNke+p+F8Edv91O8Vzj6wfIC2JZ27gXepIRrDnCWv8bcXNTC
OSnWmKQJiR2YlGMZ+rBwzV+yD5MLplYK7svM8efNyFrvrLKUp4REiN0u2k6P4pIaeWoRVL2a7PIX
eZxsrfpRwS5R61YTZknCzz8GsjSMdUYgICpyw+BdEmjhlX92j7ybDzIbxwoCYxUCaW5vxV7z77mn
ObjMFQFZHHH7mK2/KQTD2sN6+/ZVaFq3tPIrjkBJJUz4ckvmwcbFBR96t03RA3qW0ThqWqNWiOwX
et8+RMA/hI4LOrz4NqNLf1240ovASYZ5ABU2DFgnDS78s7qlIfULSVE9cNFMx3yX/Lx8ee7K9qqS
k+n22AktXXB+8boluo/pFQSEi3ipWJqmtM/jNOksiaAOxRdmp1+3VaGcN28AngIIwlOj6ZxE2Qcv
4ewJpMLenYx1zTeqU+74+J/gzF+J6FLCxHQG3E/4TIphpIDyMgMivPPmY22kGpo4hIF3Ej4YwB3f
uN/ah7Xq4mBTeyejm29Su8LcdxpTqGJ2oUwUWR4CRZXpIRZHy73GQmLXmRwVdvre0Sl86aVoSi/L
WraCy8+6xwCgrfpruptrmVJa6Bk3gBFdMIfe/O5uCzQZJeKostLsb+kc/WPkwIfcz1xQLG1Oc1g3
9DDJRcFKMc3MgYJoYG4auJPDCYUD2/UQwRhWojwXw1D0xZbK/L2x8SykOKB1CggsgDWXhkKWyFlG
gGmaa18Bh0XkoEc6Vys6aTPiTBuA+PdoSWGunHjncbSRwfpNvwqDP7QF9RPjVd36qEVOnWqIf9eP
wfwHv6kSR6vow1zd7JmTw2TlAjfjrkhzI8DCrd8L9kvD+as81C4vCxJK76y/J814rkIxJ2Wa6HyV
eANBdl/acRnT8RaQKssk04UfXV2g+bjMYcvQ4AceT0+aH0UR9ppkB+qx5lT01lz3FPs0u3CGBs3l
f49TleJ6ycQHo2cdfHqqihMiZAK/Fk0LQYeLn1+i9Z1gUZcLQ/LCRLrnR53NvEp4CCnH8HrG9V5h
O0LBNoMGjuKQfCAELw/LhMB+II5bc3Uz6+rDvn7qkiPwtYGp+CWmgho6zT/CjBWZfkan1rka2Yw6
0pFc1qL/qgUxAo8zVYqCsIi+EHTHPI+0GNia+cRlaVeEwwgYGdeVp3K4y5lTRUBy1hNpxySvBvTh
S2BiB8vZaSgAtCSEesiy9SckPs9D8egVf2mGkQ0ePpvFJPQseOshDmWmjumZXMp1A3B+s8WC0z4V
Q26swWQHHNK4q/PWOFKIpB2sPyfIRvaPYw3Ny3yzdnEvwg5RrqVyAbd37Z4e6aVLbe7hvEMuGAWs
dyfRm8+Rg/g52za+/SMPcKgMQhw1cExvjnWZSaXWQPODoCevgX31fj1u9Rh1pwp2uFmHAn09Ru4X
TySd/p7+Qcg2Tbu2OVISuMFG+vXI4fFMEiVqW6rSe2YUMDUzmcMNsuvokYmqZAeBRtU4Pe3kDEwn
c2FZGbw9m0ZbAwA1+u69cAYvtNJnDhBUoMPQmQ3TOj+8/eGE67m07vr/oUDZmqO3B4rZo/fhyOQX
9K2nWW/Ij92jDVms5FkGJUYOQAhRL1TxDOJDhswQj7OX5jlBYg9B6LpXkaEl/Md43e2iwwNKYdpx
l89D8jqnNDjmsd9dpbezmDBRRZBTsEm5W8QK+zM3HiZEZBTvF2iEe+iGWT+ciuWL4BNsCF3FoRVD
hYSP+XGu3gwfaPzpS+WGN42zVgBq53y6sV5jDsayuMBdlZqu4FfjXiDhL/r4JqJk9LAtVwbXWkeE
wGNTRrGshdarV1zAmTYYCUwOQrdGa+Bu/9MLk3hAtOmgd3YLaARuVVM3jk7Ep88WTjxJJ5WjWWrG
96xrMvfq0eb8SEJqhLgYiOWY9GGC5WO/qRV67iKsqRn+U7lobfzUBtVsbnYPIPWI0AMu4EH5ZWKU
46q3uLAXX5efGue18f3RoZc6Lw11pn3Xe2yj7GxXcR7B4GN47UpznWIPDhSthYIJYfV4s2vIkSfo
NAyLIPK9dEKNoS8fLnuqUDEV4RJRd99ZN/9r8CJPzWodkKeiYYzBK0S2o9M+lH3BV+DpYvZaRZoJ
MrllFzaGLAf9ZiEnBvJ1P871KkFao1F/VlZuiEGHLAjkYs+J1YGOhD0oZ2Rc3mZAUQdWM3mMNRcW
vzYFqVmpnHv7azrhDp9QIQ5Lp03hXJtKx5YHXpYeMqJ74Qqx6K/NGLBbqKiBnIO0Y9uIq4Gj1JZd
4WyGUjYrzXBim6wt33Z9hyfMxn6DW4XrirQLwZnlR6EZVAPJOLRzU8Evsn1MtvTrTv+9g+LDQMYf
+QyKutNuMEMFDXi7zyXToj4GND824dt7Xidbo4tuLhycR3zuHkHvhi9v3d9BQLV985AkJphpTg+F
bdxzU7G2ZYRL/aLeujn+1AEKk9yembB4wcmufxydhgJrj70/N1Agp6Ju4kjFBDFCoo5anLF8RG7i
tg8ihxmKat45hv6SwWOC1UJVAK40F1wAfnndaWRroYfR91WcAzkCPU4lCTqc7dgmVQ3HY65Vfg/A
bB0CPJe+B/1YDT9ql8jG9PCHHnLFyn05/dt1UrNisnghtjCXfEJGjxH/FLQ/ta6zaAOs8drIPzhn
gQaz6Cg/j42tGSqEehyFwaaagB3vJ2w9Xcc7pC8zKPqTZfaWSl9UsjmDk+QcmBEG+mRTpdCaaXrR
QSm2ew/zaH+HCaGh5jcsTOpRHurm92gCyc+lsTZLBhHHvA0KD03wR1A0CO7JFE8OFctuOB0VFFTH
m7bQVhK1kCBw/5s8SpGKKn2wG2SiOGSYunwDa6D0cTob9SBVpkwFQzQI+efQwoSlV/oURAERqlbo
naH+gsVXXoubhy/TsYzDeQXc62V8cw/v9qfjXItbGOBluJ5Ro+5jTfmj3Zpa2tUe9nEiRN9wxILQ
hplE/IFkxJag5RBVhuO3NuTpCxrFJ6q+8dj/bCBaJF5g9EDINVo4DqzDI9Kf5lhna5lBb8z6L0JE
q8tC41LaEtBMMtpXn2tyORqyAOMRmR71X5bIOyH8iwtyGWaoF0fBfu30WqiQfRBmt7VgLL8LIWtJ
1GhhuRTTF+J5wnatqBu7ItebNGGPf3rU1O4WEWPh1JnR4dEUkZe6aN84itxCInzkANCHyPCCjCKF
3+HZUBLnGUxL6mWyFgjd0nlUOzRUN8S8U3foG+6l0q0P4+XgXKrCsT1aAOyKsUJCJbt9t8agOjaH
01dM9HJlOzyVZC1UG3WTGH7ewL51BOC9zlf1Tvz2RILmigdSuXz22VkxbRjJwOp6ykQKuK1Yjd00
FKsfrp2Sniqao78kRxLP1lNLwCqlj4eQIYA/pL00tDalYl0iKtAOFbqzc0VnyzMiGC5xJcVCmZfC
hO/75DCDcch5Affm5IT4ugkvATU1KzwvSz1X6ewfKoNtf1o4ADyMhtkx4SvYPi8S7Q+r/pydmmhw
W7b5btg2Zn7mc1Ay+MamEam5gLqSGLomRThEopue7bmXXk7ciKeWVS8TOBUc6SIZtyYPmR49B3pL
232BTpmVlC1zRURGhyGU/YiYYpgBwgCfwSadlr/kfCqxowpK9P0Z7p1wleolhBHu8X9503bLaWPl
MeFnKgu5cyWo9pfpOq+Lx0o3+te7G739GbwXrCKi/30TURVu2VGdx7zNZBhi1uXBMx3oILL9xz/8
irn1tucSvk1gLVVF2dYj8rPo+inpH97I8M+YIY22AeKAuFg31BTP2NjBKYXZBbe905nkDJPWh9Cs
MxNmdwYg5XtzeKGe7gmcI5uUvVV96PMxTJqUK1x82MPY+4H/J6J73jS5RpmldpBDHRIhwgGSijtA
AZYRKZ2alnc0E5Tv3ZKB2EgyH4OdY1oDiyuKFQX5+T18U3zqoSPowJnGEUzbe3dEGxjlm1rQoIhT
iFWXp1x2ulU/M+ar0T7eYUueLeWp2RmsWzlE3rIf3lVGWKJXROYAFpXLt+81/EgY67pk5nTEi1Wi
CRQWuF0QfIEJjCVGTQELPf6VotJGhWxqxz9xdG+O27R9zhH3TKsrnHSGgNgOyjU4BqXLORcrJiAA
9v6/NCtuqVVtI4jE13RkfUlnAMQEIFz8HlnHTeHQnb6H8oLdGHDYa8+dml6YYtRur85pQ9/VHdea
jOi1BXSU/Wq8CvA2noRqlhlHhHokb/0KQkrcMVy9wzo+fhUBzxQMO7QcSMyWkYzsuRczdNJGVCk+
TEx2zzXgBFK6uz/Uufk2GMuq8lLnKuj/UNastfbb3hY2TJv2Ck85f3r/4MhrqKqB+8wBc8qvW/tT
wsdEjJTMC6FpyGUSADlr87P+leOWSQrLGNkX6r7VjXlcWz6uDcTc3O+p1+jTqyABEQiRog8M+VdM
4c8LzKYgAJ2YKqpNhn50j58T+hqtVCJ/giHxDuXvr+5+naoT1nj0XKoFmfeNy0jatP6Pu+97qnNo
dOc46Spte2dx4+AyCBlMldapH141oeFCcih6V0Nf+TZuROG70lyULZTo8nYQrS0nKhRC+F2CdOa1
g3j+pt3mXzlrvqf2wAxWnsPV0yageFa1+e6LyLHeP1oG72GqziGk0pGLLJCVLwAiLG5XD5XHNYZX
6PSJDY/uQI2dwVDWlZRE8WerwRcpwXRd9prDYwwl6YSST4KNoeqP8UqXAacPb86aLZQv/z7IZe7/
ddnDIuWlhyPp9oUx4ja8nCIrLYTT9gXT/TjhahFJqqJqq0F4/YgmP9c4ekdzvly/bYdPkGh9ZbF2
9iblxJouTAU9rkBeU3Qawp2D38V7pAafvFn4mkFLqlw4bbBq5lZ5J4VqJiPmpBh4SNyJo5Pg/Ig6
NMmuq648myT/kjyO49wWxOeNc0b44JUt2JmFr9+6ehje7JBjvywAnVFQuDwsG9zLlqMl65RWLsFI
q/8cgEn2DBuX+5tc6EndvoxmlGl1PeuSctQ2Twi7iHGorVixbMqvCnVDuRB0blyDLl1TnsUVunnM
SqwjW2yRcyIgXrUR3V7Nz0DzG0P+aXi3HsSsGzY5DCN3zwKMSvGYaEPnXXktMQDXjZE42m5dsf13
b2lXvdJCGwQH4HGYLyWxV7C/xu1VTnzZrWBBtOShhAtMAO47fPlPuJtPb/xf/kOGblvg4GWuoymL
J4Od//ultVh8rd6F34OstIjuQavcUts528yYlUYirlvjHjb157lJCvrrnc670ihXRmouRXGo+6xV
b2S+WGrye6RvkIktRkk2sN+FuUht/pDSzx5Mi5LWQJVLNskm0/6+vgXfFfq3lVYq59YICwxzm/+W
0wHvBSrWtSSFSPpcjDYyVq/kDYFj9uYFNHKZHTIZU6B2wuTTpRmQZX399Xj3pG2UMHhUIRCleBKU
sVuM77klkBLiP1uJ0o8hnQl7TxOjrqDumqXMoFNEfUhlRYpKq0L/8IriORq1VCkrhLknYtnNtsdN
GH0t0biYtwSNt8QqoKaw+ORmDOrYTDG7tw2oaiTYBQHJfkKgcuCVqI2hYufu1mX6m0J3sq5opKRt
NOorNlL8ho4p2KDVm2qmKbQnWwGQYeiZPPnI1TdNH+o/bWf0+RZL4QCDa1YJwQGLBp/O12xVkjZX
OxpmDi6S9j6qn6+I2Ey0IH2nGyMQy3fJ0A2rc4qCrLvgzJmkZSVldofZaZzRuVMuv96BSHhXNA1G
fluEX7xmAM3YBILwh3b5jgW6IbHmpPjM2lNyjBy3TgWpzaLLS3HkjcFKWyFxj39vVjJnAyMkMyRq
VJlYTCCkB+nCdcZKbKX4p54TtyHJkwFPSWgetQnDgSti3lU8GWU0bPg2UQPdoYgcEkrThALBp5GR
skE8cepXj8wuJ0ScFMitTetTvPQEuinHoOQdj7n7dKDpLEqjAdtjUNGUkrvHs1+MB/k+bXkkik/O
cPDu+KEt2Qp9ZdIBITRv7Lh29pmNqhH05oL1T97xJfxMx2kejf25y4jyolz+qjUwKyZC36+SllmC
Zb3TkjxFj+0Lu8m3ykV+6v1ezd6bjKKYLGsUMZp+8ocxt6nerV8dsUw0GQtNT0zfUjObsVJ1bylR
gNQcztKC3/gorwUymK1GL4drgyiU4prwci3R3KPXGNEIZsu+xzzw5v23egiDtfdla1FqdFsA0bdn
uftUc5iPtXdN7BdrdpsT9YCHuNll27aw3cxrBe/uUwI42uCJdcpV0PoLtA+RpMamYg8XVoAgHxRQ
HFd9yU86YQ633mnk5Ueird1ARdfps9MneWb1aouaMh3l867CFnm3cMH1KhweFN+c36YESdofLwgO
MoM2Syi5t9wMBj+hh+k6ioRIt3CPLmt7iblZ0b+EFdJs0jZGWB2I5K1YSddmshZYtP5G1rMI0tDN
mW9wdvwb/Af0qK4wYJmu96QVeEPBvSJfqC6Cy3PV1I5m8tT38ghMfVDv4/1GaRSa3e/tkY9A0uZV
xum0zdsbe2wE9QLzc9uEV6dtpsyWW4iFkOv+zFPwO4kjmHtqt3v5XjxXldLgasWAeHWHRxMMLZJw
zgb1zGp1u6s7ltyP6RhLUfvI8y5Uw3fo1HZXOMIJgGL7vz0oSUJEsFtNt4I+w7AKxBt3RRBQaG4t
LZh666majEmNQJcziLKNVIaWlfYsyDzLEMDoiC6fauWoNlbnauHO8u6IAVFzpyxonw8QhXGMZyqF
YnyoCDmtvlw+9YAsMPQxG+XKhI81gzczHnnneR0NhpvmwCL2ySQi4WVcyjfHeFxZDwUu4HO2VJA/
WKw37IsZ2PwsrtKV8i+VgUANJAGLQgxtOu1SVIPgUUttiuLApNmSFwmIemsjzRgk6NLm1XMtB/83
JC+i89ygODN0DIq07AGLTbDE6U3jUrFqDGe0musqhTda0notNTIsPwULHSlUPHt2IBhrsxPFGMEv
yuPkLHuE96As+3XzSB/3WICYbRaPOtEfj1o9qhPUDLXGu6BUJ4UjCq6P2+oxIM49OROyAxMHBiZ1
5Lkq+Hp6ZDvosETxUFNNxafR0nFeZ80SgJi7Y5HNQ8X7eG0t7m4/8Ewx2UUdpCciE/iSL9XT+WGk
LCIIZ8R8HOqo8IxT+B/CbcpNmAEDYIOYPnwLQmYaavWjsZCgB6XcGR0XUIm7sWPe10pM5g1ft7Un
1nlAqOgu+ptWk43qppjhtrfLrl7qJTr/VL6lAZ7sJSU1F+q7USuXirr+uBqUtpB+cm9MSTE07/mN
65Zad8v8cOJTQv/ZSL5UiU8XHsqEWpcGgIYWeR7m6hXW/LjAQKRGBpDcHcuwhc1NTB16vLQhUMud
9IRJQYITfSdn4Y/+psMTPQQFxpIvVXK94XUhkdBLQBw85DqUnrpVZfF6zq8o9IrWV13u9UFnPrps
hKYg1mhPfFKcmWSYUiCjJiOKRFlgZ4HaC/kM6jNFGX9YHaDMxLjErEfNoENcS4nkTS9WpII0eWbl
oPR2+vLS6pitiiLKGYeWnd9WMI8fSEL92RhwCoHbswGUsXeyiUZWlri08GTXPGHIItr4qlFI1ubc
HBon/SXldYgz9Rzkr1wrbZ36qh1UG6JYn5bSy1Obg/m2azxL4Z/lB/ely1ycFcrgzTw36IPx9lqH
sWtfMT+ze1i4RQXyJnQsqZOGBo9+c9QaG7233r1+8D3aZOfvgtc0L+3Rwi+ss67AcZzN+zUHCgj1
k2Za2491iTh0tsHL/Z2pUF+b4Z0wanjf1GXjpxFJyzVl4uoBfOpG7zAmQWi4w9kr0j3fd2l58dQ8
fW9fR5R7pVsHbcdAIlPPA+j8mpXh+j3YhKTPnL8+H3XXUAChQ2FO4uyVVO2bG/BDRCk3VxEZsKgD
wT49xg4m/nF54Xg2Psr4nch1j/gmmaUuAYh0wBezO52iEEMGPzF+Zc0NI52RTyeLV818uAB4prnP
wTON+g4yBXF1BnEnvVXp7VcdXUsxbRy3M4kiqr/Lc+HFByF50yGYkMchBWyZIGRL1zcp7Bg+3zEn
NZmWzwRYD3yivY4fwjLqe2YJMkR0kEoB0wIX3rD6lqspNEp1YNKPkfQhqv0PbaDr84UKiuHrDBmK
ZG2RvS/Ofwks/DXaCvgbm/vGINAQTnN/RB/hu3HxbS4INeXi+n7RYZvjSuPJDwQtg6uZOeiE/k3/
pFInNk50o6shWrTtzx6RB24l+DiXckVfLaOlMP6S0xLaw2J5aLbXHWfUGK0QBBXcqPziteim95+a
nJiZS4j7Z/6UPZbK7Rr0O2niC/b627bbPdOzu6DULbWtJNRrIdfSGODU/5ZQhMEY1SiPLmPEQDuh
TN8aioN8VKzSrrBiHzDX4+wBwwovFqjqFQJBigw3F7CMdHdrygOrDZc4sxjt7kxaPjN6wMxYlokB
ekHPgPcAyhZ58iLdgRM4r/wEqhWyr5vn+Wy7y4JTtzn8c629bJ6nyxxrUBxszgnA5u4Cro36adOC
wQcY4pV/hyjTLuUZhcYDFQIJwfxGeNxhqMNxAxzpH0aFSPOu3Rxu7Gk64WwKWhXx/xLTIu//2mxx
0gTknzrvmbAD9QHQOU1A1pGDitheJc7g5Bq7pN5hTuBwUzcHCPTECPOURGVlZktlUf8xWtMGUngg
0gyS8m+AaJm7HE40I+SiCgLmv5Dl7lc236lk75mRHxKIAMEXOWd5K0PSE4bmOD5yqHyCVNR3txwC
LFPdt9a75v1sQgHt1ugJNU1dsu1k7JVt00A/ono1rlfgxB3WXF/YF3X70cBT5ivay9HWBoUqFY5n
mLOVljWErcoX2s2KcrTPjKE2YrZhNSUxhr4cu1297y3v8zRwsjU4+JH3bkeE9BeHNRAH/e1ojhnm
Lo2TKAdM8KmlqSiXk+jEMf+3WVpzPTAjNETT3GC23sSHkUfQ/Sd8UNTVgFuQLhOedM+gRhmiFZbU
+iBhC9kKVJZhoTyIRyFhGF8sMN0Vg1DkrvBWSd1HVp85+EFMDzFR3+V93Dx1dYefgT1uyhfAPIVP
lsl1tvzG5I/hLfHWEwJqWicZwWZvMxKosjJf3g8i147yyLo9GB0hSqnjbM3V3fepThAuKTdG9o3N
+8jVt+1OHV/T+JlPAuYrBPyzR7bhb7LYjbm9tQ/ld/FL6CQwJ6jwrPmPKOX2je5X25IqQ6S8fTLx
C1XlPRAnz4yjmBTeK6tMmH11zy10IkLP0WRZbMSMSIrtKhxCaVLg4sqeoQBA+RCuyd5At+FvHeT0
WexTHNF4MzKnLbAAZYmJKw4djJn4dhPNF7pTj2w+Y1J7Ji0MAY86aiuCY7Ym8U7vvBett2qNv6ix
SBtgaoGh8Jt5yMN/QESgkcucvTxkQNqVJHn+ndO/Czkokcb+E52LhdaJN8R76+0E7dr7CeuUgFy1
gIET1bASQb/Jye37IMtKo8hUGooftQ6hgUjdoe2rPOKaAdLpI92M6JYy+tfH3ejzG0AxAcIoot68
vzdrk1mSzaOLqn26KHlWhX8fscgfd9Fyr3AYuTVjWTgf25uJnvxJNcKU3fGCO208wC0x3JcQ799B
VIP68oHnxk/RjWHwiTdzyKGvoIZup7VjsdRjBs+Glp2sXIe9OFi7SQMBMtsUTGkHLzzHHP/1F40L
v4uMLPsevwfBGR0N8k1RSFtS3TsJQJQuX78605fD92WeOGVTAHQiQH5Oe5H4VlYrscHvLdpDbEjQ
2On7DXhmmPNll0VszfE9tEgrorCUs9TOrsXP1EaSeCnxBejrgcLm1n1Wi4WIAZmBryq6O9u5HHNM
JP/q/Ya22G7sL/VndScbbTNXp/v4QytlLu1MGDFBhpUh8RVQTLQkusrvDMwv0Mj9PjkxgPn6CnjR
zaB9vLOEkmUpU8LGdXlguz3wSIRv1aMYo2iWAOy5/qoq1e7sR27Ssf3FZ/WKC5PXYeW2wW/sgy5s
+Xc7kDbxJEHNurWUDxEbyOPskNlKFMpg1vlgVcRzbdhz4W/HGI26nmH/+qljzB/GOzu5itzP7w6H
ekVa2qJumdQ7JDsCLX7GIFDcRLyojBcWxD9o0HduITdIi7cRuSal3YPLI/mBFZdgELhWWsEZvE+C
KEq6WEMMYaydYs+CHFK03sfaMA1QYYLTYHDW4M2eFilSRTw/fo6muIwScXzPFyxDa3Ono0BieJ0a
4EbFZl2pckW52qnrZpnXRcKQY4Z4PftLQwgRQH92RnLWciGtXaI6UgLPwywPo+ad82f+KVmT33RR
a8EqYv3vISEwwmI3dBaW/+4FJKn4izis1+aQzQf6uX4Xh0wFjmUQR6KC1Owaf2tKfC7B0Dt7bHx8
k117o0xjNjEhinzAV2qfussF3Z28bLNBLV6kxw04j2CG6Y+5dLem85vdIjurOoso1YEmKSglxcfR
ezjhd8JA71rsAVjHJmmjfB8+SDcirYsegAhNrTqiFJvu3N5IMHRAaSxTKe+HFBuuCKqU1EyiZPlc
lGnpobB006MOMDJRqm6D6lAl9yUmSLyCgBW0lnfMebdd/5UkPMXZMnUQCZM4Xw//fY4ixCom6Ab3
ZiHSP+wTVOzJbi+b6ClMMlRu7sif5vwSx9n0WdW9Is7802WIlRbS8vPqPI4n5gyEbTFNat3fMhOE
FGKVRdlJXShoibUd5YOO3MjmJi96NACyUtGiXL83FEdboNSX40n+tp7TdDkTuNmVyM70TuNg++67
qF007QhfBAcEbDWC0YyMIXgM3z7dlkLio2HJCr5e47x8vXeypDZgimLfLJ/9MecVQynWOWKiGZoR
vETT7KLRxMX/45H2dIDsFgRMnsMz3C2jfwYoiQnm7g67rT7Io7V3+oa1Wnh1eBHjRig17A9pv1ED
3PNlnQKjymVwxSitjuAFS83VblFiaFhcuv8z36oEjePJhlnA1bXV6ffZo8smsS/KDmeCKvcsO0F0
59YX8vN/oMymnRhKe8sjF86T5+nE1fG+BJBn73wPmuHcS1c1A8xvfDSP0QU6IQk9EYIjPLJdIm9e
CNEgMGm3+rV7PNUUphG3NHRcAlHnRBhj5tO+B10xf6Dcx1nKBSKJ248pqmoxBb/IFo95PrLL8kb7
SBg/ey/k09baFXnaL+WPfHPDsiXfyjZPhY+cC2fESY8Fc/0qPKh19k8mC1xZYlaFkU6PvTkIk/FG
iLSIXiqPmrJbEbwxWpdSNBxjOGDtRXUduxsMpAQVkTM3/OObKI7ikttTysxlVHPstSJqg+5OvJhw
k6mbLwU4iTTO1Er9SonUC7LnZPFXiauHXn1yWR0QTteu6WiiPuiDrz7K+1DqAeFNfPE5Xg+uBh6T
WGUv4M891W3txGtweAUbChRwKSbW2SuSrvGMK8rZwY2IG2b/RnTEAt0b53Yl6YfItN7LAgMHMg1d
qD+bES4Lq4e9wzv3Uj2t25xNA2NGnvFOMJ3IXbJH/k80MEFKN6EdIWUC2Y9RsFrBOejMT1JzV2y1
nOPsXELVSewlnmRgS0OExDAOixtN/MliBM9hDi6Cn4ms/k2P/NgIyySmEbdNwcEefoh7afXmUwBS
1Yt0WTQprY72J0IR+iiywf9BPaFcSGRQlJY3bQv79RgJ5yPrPDmMG7N5jfGyQUqeRgzRz421d4WY
9bHQKCD7ezCsEf8WmmVXCLhDvJEzU4nhxEcx9e0sq8MUoVnG+fK7eucgEzi5g+P/ZIhkd33RggQB
TqDDsnWBMIUdVXel7g3UmiF7t5LFk29Fk9DQUdyhrY4Lfqt3ZUVmrLAZQUwmu/St5Q5nB5xJJF0F
rfz9JjfjghuTR1kcNtxyjZuKEAruyS1IygJXzMiyL/CEKd/w7cPiwROrmdvFbrgXGI6LdkBh6s9Y
FJQ04NfB2gWb0YlnEOW7x6nKX9vCR+7Y/hUBwYhf+jFRMrhspms8GVcLxyewRJPjHWN3EEOWFpuE
KwP+fsBx2PW7ywa5k7mbOFi7UCSGZKXUsrZWrATRaI+mOp2F58nTHfMDZiq3qT90Xe4M5K6GziSB
QQByRugIaUoCfClOO+YwlpaY99ZMTOILIWzlzy5AVkOlubxvR6AzebeJ95UhQAboETTfrN9ZSt/1
FtEuyli97BIdBz3F2TYwWjaZkX5SdoJB30moA6WRsqIwnqHAQ28iHbRqSR1RaDaj7ON7jNH9qgYK
U70erF83NOxyzVRqtR+W/CoMBLlzGfSH07I1kIKw3KQN1QM37naJFLv02ACIWcu5lMQkDgcL4gFQ
pmZcp16Bs5ixlAnWwoI3IZHC/LdlfThiDovrlw5TnF7nGZzBjNBw0bQb6NLVwxH0pjxz5hdz93wL
Ck9p9T0HCzxl9w5PB7rldHpnNeNdisiMcgsZjv922VVTJCNFB63hyrkftZAV3/QYWLzR2D85yRyY
zo8uZf5f6mnvU+zxETon4II67zy2SimnVukrGHPFEsrMxCWfenUM6RT+gtYiKX0/E7v1KZiIUEwX
Q6xm+XXmrDgB4wW5HmUXEXVS6b+aMj+cIgnR39C0PHrYSuRfvWcGRIYJ0JikeK+z1RxVHu5DMTCH
ZJ7MM5If3DdFD//Z2MwZjoSXGWNpxAcqmvTM6/KIGfpnU/pY6HXtUOj/AQyasoDO+H4tKusdnjwv
vEKzXya096fy6s1fEY4w4zcHNjBFfzbvSyijEZn4Mkolp3OZvWBZTwykrVWmy4iWCsiFToCYtl+L
TfZmvK+AQHRyDqn2YkUtwRjBwieXkNUa0JOC7Eli1IBe+wFZQwUnX5obdoazzKmh1UC4SEGCYh7i
ZUKlMHKgPy85cdpLaiCp2H0oMqhLNmDOi2dn2IdIhSFPrqWDuZf87Up7i6qIS3Rf1ZYX/0zokXJF
Teu8UHllDkIUYtYkV1GmnH3xAIowSmspHQBeJG4bsvGxGaIQfeghewi1lyVqCGtyvETlCe6J91zZ
1BJ9rK0T4u3w1ae7aNM/IqpnKXuHnUkNO0dRUIZEgaK6xObn8BhO31n0oNCoQ166Y2AM8lklO0jw
6mljt8Ey1ftTw4d4lm/6+icZdxmquxo5/mzTBMDqXSeZfudcuMjaL1rVoZrGCpCfzR6eyiFkCcRZ
i66vjHV3fuhHwVgxU0ES+Y5nNYCH7DxlCi04yVhsmulQGoS+RRloCB14Nkf0xEO9XDUVLp3Uyh5B
WAKi4S7HneNDRJeY3BITdPdXb6ucXPu32vUzHDJHEPkWI/HpcptTqcQhhZKAgimaFni+0h7eyOku
UyuDm6b1i5W81xkSVaMV3OSgonDpv5MEOhpZE8DPZ32O9NXFZQv6HVuFiSRbpbVMlDSSoptUIdOi
bAzolwzll0PXHDktXyV4ZmSJBQ8WQv3VBWdp4t6u43YqU8fXhgMQZlrdqqBKxUmE7J0zALqHexln
HD2oLZlrLlFvx908e1NGe+ssbo1c+mYlC3Jo1Rx+0A3qQm+gy0uU8xMW+SajT4wkmbqSoMqWUMno
Ill12g/BqN6wSImml/G6qEqbi98hjbjYPfFLW7KXOqbgx/iia33e2dQ1z9KQ3P64D3PxiJgqcIqm
yYY6aog7sXT/Cm/Xf/+OAyAMlyzavaSmLK1SJa/9+4bjH1ahpPlxDd73sggNWwIr+q2Ta86bEyaq
W/M8tymiAxiv6vWQ2a6QjgyRH5zLMpx81y50zKN99M3rBlZc2qFAaKnJJ6+DzqRlE/lMHVIIyacJ
b3Vjn69KVTj8S5CeDRoR94R4xv9ZqzGy3Oj2Hh+aGVv8RWEjpFFylwjvfBWQbQgxHno/FGufLlns
FWFABRvjSoVjIFsL2Gpcf6gkT0k2EnUBgsfjdS1aTQwg0B37msm/CE/Ymr9NPXAbCS6xPAy208Pg
3Q+uMcQk8OEPL+1Lrp7Aus3b4SVX8t+PDRdQTppvU178pu9zN3ZjRL98yOOX84ni5BxMm1NSwKRI
4pfmzkijex9QRxFNZBZoCE2xDQSC5yQ7xMo/fVFhW0Iy5qzFAHHSxkTGJCRG+gR/8TqBtWmP7a5U
BbqMQlb5FgNEz9eXqTwxrSOeZM6rlP7Dexof9jIAZru37cDg95cBQvNaJ8PukHwl6ikYmL6Z5z+S
/QJjfFom5DZxCOqeUpcYBHH4lMzf6uX8ARbzwuLc02wEg/Lb9Nmigg93+ZzDE4Qjr94Azj3gZKHd
kTBM0sKj2voR+PNBmPQ7OB8BhlPg/BPw1g7hBAjzyCLNbjfLCaDRT8DrOuwPJGN66hI21sNN15Am
xap3hb1MpJXI4Kr0+VhbqmZ1S7lp52baFm8pPsVw1Qx3EOqrIRqDIEgODfIlMImipPpO43qocY9w
FADP8ooEbib+FwxYiajkHLgaa4/SlEBVABLbwLoCUs+ahgeJYMQZJyhZy6BO92YUzoX63WCwgeDn
YYn9DAka7RmKNDY7irPH+VTMbpwQ0ZTYeGvlWIG13v/EVU9uYIKLx9o9arDghbiJAoo94GCHDU7x
y/jGtU2bydBT9MIdX5eYlHz/MCCPhXquNnQkfiAfU4xnFlY8SiHEfCv6gKw4tvWqikgvuqkdsYEY
TkW70MKcRHwWX0GCzCMaXeVKRw1wZfGrPhjihnkScRT8YV9zaED9Hi83LRKj9P1J1wlAQfHVLjzt
uBv0RgaaXy4bFUWYZWkpbKntkOqbVifSorzb2TQhMybbuUlKcm4YkrNlK59YKLz1F0InjtEmvOBZ
cDKlkFEPGEvOP5Rqm1OUNO2U5pCZ48lOIcm6PqO97GfaZEsaKvVMIApTdYaB6AGtFj1RzZGjQplZ
b5M9Iqkw/M1v5BRX9En+zsb2kUWnWa5M7fAiG2bTLR2NLafR2zIZMQjmwa3TvCyvAk3DYt7YYZo7
5Ly4B86lst5+dXfl8kz3iyK3Dj8Lgl36pZYZeRcLs7Hlox/co1cr4CCaFcpOh0t2vRyIl8n0YBWo
nbyELuyh5L1vIP+K0KPg6rF4F8w09CkYT2E2JyF54ZdZ9QpsL7tBevAwEW5NM6cdS42YXmm9yJG3
f+dCS6kMAOz8iW2tTnlHZ2ocUTW/Jw4csNaP/hW6fO7lwgOFdMk2mTjMS5eHFzU0m8tsOdh+LKam
QB8IgiyYwRW5cneutFCQ5uOyWlDXnSarSzmhuTQRLkY/flcGIjcjw1ylML4sbw3JDa7oReDzk0oG
+cJ84iHLgmAuqRRp/xhM1dv8Glh88eOStfLNMNw/XkkyoVfBonOLFj4w/DGcpPMVX5I7Z6X+ESJ2
UqVVXUSaUaoQGwr+VNL5z0umvVhJjow/o4uCojtInYVTLn72VH4GnxWX7jIbeL1etFsNSahy9emi
yW+AtaYgMssUN3oA4HiEjoFWpoMENxpUomBRvwoFj6uL+cWFxL9XCi0Zdhjj86+WDon9dj3+/xW4
30bS6/J+h1I70nJfOTHKwucEMSQkfQCtxxPf+g6cTra7U+237j71yKTq4YSzwKwsVLV42J8xu657
DWqjvKkv/+TeQ9xtY8Nz0JCjXDFJX1pwVRwwwA+Kxg2UUW3UeQLUkewU1LTRznB7Z4oC4WBei2kB
RFLXxiy/IpWJEQJBJUqH5NkNrouW7Dzg6G5nw5CF/2+zXkVU820gnZnBfWub6e3hCnozwj7zYXhj
XfQk33JswEQw11F0HnYMDsLUeck78zQYaL1GmyeFyU5Ts8fFVxXe3Uo1WUvSA3cav8n5RorG83Fm
jLIAEPfRTkcAZO8qlBm3F34KmNA4RrzMG8wVQJsvCX07ZiocmQhCnHPle9/HYiR1bX85hela7MGi
/CfDq3ZX4zR3rzspBAvBp+LlOqGQIviluFcMmUww0sN1K4M5gOJmKjWymrCvWwBarY9sxFiboUms
JxTZB4XqEb6EaYGTJ8mgcmO9f3Lc5PZ7EjAYRwza1geV5SiNmIVbaLAdigYxOYQyOfoVXRKoH7iZ
9VWKSE6fc2+UTXxJmeP2Ivm0+oV6Fp8/AURDZlvPlugPlFHoIksYKycQJ3QDLTOjD7Ed+v8lHavQ
tzHMZKedGIvJ9Xj+9Xp6mN11EXlOetBDn8+zLzam6He6HDEn0GZ+PJS4z6RzrWmc7wA/ZbVQhdcN
11BkT471RJX9qFAQ6ilVjt55N2ldpl/Jr6/8SJTQilQiNWZJFqttfXdjxqtz9PZ7t8uWi5X6r5rO
9P6otsH8LHHOSE2+dIYf70gvn0RMKcw4NrrmtQyQErjkosMbmVsKPqidPczVl5DGtpMnS7J7qxGq
GsgEH+qzo1OS1RvdF+XC0x/acfio/rQIPxRCL25kjBNV0DIC6tdk+sEFkP4t+50t7Xzq7hKhLNWq
bF+UR5qKrLPu4VP9exx845xHwhLt6m51cnWuwVl8YI/hZCQ0yTV1CCjoX8cbSsS18QAeKpdDu8MU
Hibq0Qak13rRF056OjlyO9oUQdg9H/KngnGUxT0cEMvvCaocUYEDoKyv6G6zv3hrgWOUO3ugloZJ
jbu67mO/fE3bsb9nSHMKzV4K5c1tLjmjomscAwoAKD7iT/ZC0HGNhMaBWP29eihPCKpu76Aw78qy
ThsxPoRt8EnXCelencxa2sCLniJTw1edH9xDJDbbUIjb4Dm2OhMsb9BUzY8Qsna9ZlEi03SqDl2x
IYKdJKfMCyicIqBm/XVpI61nQ7Pd4PoNllSTMXzUplN9vX7IgeJn9Ko/jHKZbB6ZPzLKmpN5AgNS
grKZspXLCYokz0kSW16UQ1NLEMkJ+kwQcpSWeGRiJf8tfosHaxM0nw/gybES+KiQ//ACAeCcYD7T
/zDMGyoHymJGI7aDolQHeJmXr0AotCP8ufWkWY5k+McCJqOLKMDahPZ2hFhYTTE8eAfpJCxNajLL
4Lv343mEStLUr3XebvY52O+fY7S51Gm0mE3voPYqPRIy5RvbLyHUxIoxWVqxjCFTSyBkh9GFRQqC
CUqR6Gqx+zU67UOWeeYaoP6V5F8Qhxnpg15c0vj2n/B+Au+spurD9Lwl+Ly+ZV4m33EEM7okr68U
aRcFNWy+Rr6GxiJZYySEtCpIGLMzX92kuOm/5lZghb+KzGXMd/RMwHSY1uR+pmjdvoEIGipT1osZ
aEpyeJwBocSc8+bP3tIjGMoxSxlqM5lFHL0kKWJgLHO0Z+cryAEAo81qvdLWxvWYGfjGvlJuGlNs
KBhquhxTF7OObxr55KgBUi0Je9FfdbLhW20+EVZXfuSQv1nYpVEOlrcjCk7kLdMMIvj7ePLUnh6M
T+Y80RkKjEKqiP75pqqsbsnsS08fbC3mnctL9yjiuEOizCdvY85A2Acl7qIYJr6YEcPd9IpMFLtG
eVTAXmufFrhEWZmFhkGjg9z1ECKTii/3J47RzTHzWQdvtYajpQ==
`protect end_protected
